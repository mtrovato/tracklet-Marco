
`timescale 1ns / 1ps
`include "constants.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 09/28/2014 11:01:39 AM
// Design Name:
// Module Name: Tracklet_processingD5
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module Tracklet_processingD5(
input clk,
input reset,
input en_proc,
// programming interface
// inputs
input wire io_clk,                    // programming clock
input wire io_sel,                    // this module has been selected for an I/O operation
input wire io_sync,
// start the I/O operation
input wire [15:0] io_addr,        // slave address, memory or register. Top 12 bits already consumed.
input wire io_rd_en,                // this is a read operation
input wire io_wr_en,                // this is a write operation
input wire [31:0] io_wr_data,    // data to write for write operations
// outputs
output wire [31:0] io_rd_data,    // data returned for read operations
output wire io_rd_ack,                // 'read' data from this module is ready
//clocks
input wire [2:0] BX,
input wire first_clk,
input wire not_first_clk,
// inputs
input [31:0] input_link1_reg1,
input [31:0] input_link1_reg2,
input [31:0] input_link2_reg1,
input [31:0] input_link2_reg2,
input [31:0] input_link3_reg1,
input [31:0] input_link3_reg2,
input [31:0] input_link4_reg1,
input [31:0] input_link4_reg2,
input [31:0] input_link5_reg1,
input [31:0] input_link5_reg2,
input [31:0] input_link6_reg1,
input [31:0] input_link6_reg2,
// outputs
input [15:0] BRAM_OUTPUT_addr, // 1 for now, add more later
input BRAM_OUTPUT_clk,
input [31:0] BRAM_OUTPUT_din,
output [31:0] BRAM_OUTPUT_dout,
input BRAM_OUTPUT_en,
input BRAM_OUTPUT_rst,
input [3:0] BRAM_OUTPUT_we,
// Projections L3F3F5
output wire [54:0] PT_L3F3F5_Plus_To_DataStream,
output wire PT_L3F3F5_Plus_To_DataStream_en,
output wire [54:0] PT_L3F3F5_Minus_To_DataStream,
output wire PT_L3F3F5_Minus_To_DataStream_en,
input wire [54:0] PT_L3F3F5_Plus_From_DataStream,
input wire PT_L3F3F5_Plus_From_DataStream_en,
input wire [54:0] PT_L3F3F5_Minus_From_DataStream,
input wire PT_L3F3F5_Minus_From_DataStream_en,
// Projections L2L4F2
output wire [54:0] PT_L2L4F2_Plus_To_DataStream,
output wire PT_L2L4F2_Plus_To_DataStream_en,
output wire [54:0] PT_L2L4F2_Minus_To_DataStream,
output wire PT_L2L4F2_Minus_To_DataStream_en,
input wire [54:0] PT_L2L4F2_Plus_From_DataStream,
input wire PT_L2L4F2_Plus_From_DataStream_en,
input wire [54:0] PT_L2L4F2_Minus_From_DataStream,
input wire PT_L2L4F2_Minus_From_DataStream_en,
// Projections F1L5
output wire [54:0] PT_F1L5_Plus_To_DataStream,
output wire PT_F1L5_Plus_To_DataStream_en,
output wire [54:0] PT_F1L5_Minus_To_DataStream,
output wire PT_F1L5_Minus_To_DataStream_en,
input wire [54:0] PT_F1L5_Plus_From_DataStream,
input wire PT_F1L5_Plus_From_DataStream_en,
input wire [54:0] PT_F1L5_Minus_From_DataStream,
input wire PT_F1L5_Minus_From_DataStream_en,
// Projections L1L6F4
output wire [54:0] PT_L1L6F4_Plus_To_DataStream,
output wire PT_L1L6F4_Plus_To_DataStream_en,
output wire [54:0] PT_L1L6F4_Minus_To_DataStream,
output wire PT_L1L6F4_Minus_To_DataStream_en,
input wire [54:0] PT_L1L6F4_Plus_From_DataStream,
input wire PT_L1L6F4_Plus_From_DataStream_en,
input wire [54:0] PT_L1L6F4_Minus_From_DataStream,
input wire PT_L1L6F4_Minus_From_DataStream_en,
// Matches Disk
output wire [44:0] MT_FDSK_Minus_To_DataStream,
output wire MT_FDSK_Minus_To_DataStream_en,
output wire [44:0] MT_FDSK_Plus_To_DataStream,
output wire MT_FDSK_Plus_To_DataStream_en,
input wire [44:0] MT_FDSK_Plus_From_DataStream,
input wire MT_FDSK_Plus_From_DataStream_en,
input wire [44:0] MT_FDSK_Minus_From_DataStream,
input wire MT_FDSK_Minus_From_DataStream_en,
// Matches Layer
output wire [44:0] MT_Layer_Plus_To_DataStream,
output wire MT_Layer_Plus_To_DataStream_en,
output wire [44:0] MT_Layer_Minus_To_DataStream,
output wire MT_Layer_Minus_To_DataStream_en,
input wire [44:0] MT_Layer_Plus_From_DataStream,
input wire MT_Layer_Plus_From_DataStream_en,
input wire [44:0] MT_Layer_Minus_From_DataStream,
input wire MT_Layer_Minus_From_DataStream_en,
// Track Fits
output wire [125:0] CT_L1L2_DataStream,
output wire [125:0] CT_L3L4_DataStream,
output wire [125:0] CT_L5L6_DataStream,
output wire [125:0] CT_F1F2_DataStream,
output wire [125:0] CT_F3F4_DataStream,
output wire [125:0] CT_F1L1_DataStream

);

// Address bits "io_addr[31:30] = 2'b01" are consumed when selecting 'slave6'
// Address bits "io_addr[29:28] = 2'b01" are consumed when selecting 'tracklet_processing'
wire InputLink_R1Link1_io_sel, TPars_L1L2_io_sel;
wire InputLink_R1Link2_io_sel, TPars_L3L4_io_sel;
wire InputLink_R1Link3_io_sel, TPars_L5L6_io_sel;
wire io_sel_R3_io_block;
assign InputLink_R1Link1_io_sel = io_sel && (io_addr[13:10] == 4'b0001);
assign InputLink_R1Link2_io_sel = io_sel && (io_addr[13:10] == 4'b0010);
assign InputLink_R1Link3_io_sel = io_sel && (io_addr[13:10] == 4'b0011);
assign TPars_L1L2_io_sel  = io_sel && (io_addr[13:10] == 4'b0100);
assign TPars_L3L4_io_sel  = io_sel && (io_addr[13:10] == 4'b0101);
assign TPars_L5L6_io_sel  = io_sel && (io_addr[13:10] == 4'b0110);
assign io_sel_R3_io_block = io_sel && (io_addr[13:10] == 4'b1000);
// data busses for readback
wire [31:0] InputLink_R1Link1_io_rd_data, TPars_L1L2_io_rd_data;
wire [31:0] InputLink_R1Link2_io_rd_data, TPars_L3L4_io_rd_data;
wire [31:0] InputLink_R1Link3_io_rd_data, TPars_L5L6_io_rd_data;

wire IL1_D3_LR1_D3_empty;
wire IL2_D3_LR2_D3_empty;
wire IL3_D3_LR3_D3_empty;

reg [5:0] clk_cnt;

//wire enable_gen;
//enable_generator en_gen(
//.clk(clk),
//.in( (~IL1_D3_LR1_D3_empty | ~IL2_D3_LR2_D3_empty | ~IL3_D3_LR3_D3_empty) & bc0_i ),
//.out(enable_gen)
//);

initial
clk_cnt = 6'b0;
always @(posedge clk) begin
if(en_proc)
clk_cnt <= clk_cnt + 1'b1;
else begin
clk_cnt <= 6'b0;
end
if(clk_cnt == (`tmux - 1'b1))
clk_cnt <= 6'b0;
end

wire [1:0] IL1_D3_start;
wire [1:0] IL2_D3_start;
wire [1:0] IL3_D3_start;
wire [1:0] IL1_D4_start;
wire [1:0] IL2_D4_start;
wire [1:0] IL3_D4_start;
wire [1:0] IL1_D5_start;
wire [1:0] IL2_D5_start;
wire [1:0] IL3_D5_start;
wire [1:0] IL1_D6_start;
wire [1:0] IL2_D6_start;
wire [1:0] IL3_D6_start;

assign IL1_D3_start[1] = reset;    // use the top bit of start as reset
assign IL1_D3_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL2_D3_start[1] = reset;    // use the top bit of start as reset
assign IL2_D3_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL3_D3_start[1] = reset;    // use the top bit of start as reset
assign IL3_D3_start[0] = (clk_cnt == 6'd0 && en_proc);

assign IL1_D4_start[1] = reset;    // use the top bit of start as reset
assign IL1_D4_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL2_D4_start[1] = reset;    // use the top bit of start as reset
assign IL2_D4_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL3_D4_start[1] = reset;    // use the top bit of start as reset
assign IL3_D4_start[0] = (clk_cnt == 6'd0 && en_proc);

assign IL1_D5_start[1] = reset;    // use the top bit of start as reset
assign IL1_D5_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL2_D5_start[1] = reset;    // use the top bit of start as reset
assign IL2_D5_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL3_D5_start[1] = reset;    // use the top bit of start as reset
assign IL3_D5_start[0] = (clk_cnt == 6'd0 && en_proc);

assign IL1_D6_start[1] = reset;    // use the top bit of start as reset
assign IL1_D6_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL2_D6_start[1] = reset;    // use the top bit of start as reset
assign IL2_D6_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL3_D6_start[1] = reset;    // use the top bit of start as reset
assign IL3_D6_start[0] = (clk_cnt == 6'd0 && en_proc);


wire [1:0] VMS_F2D5PHI3X1n2_start;
wire [1:0] TE_F1D5PHI4X1_F2D5PHI3X2_start;
wire [1:0] SD1_F3D5_start;
wire [1:0] PT_L3F3F5_Minus_start;
wire [1:0] VMPROJ_F1F2_F5D5PHI3X1_start;
wire [1:0] TPROJ_ToPlus_F3D5F4D5_F1_start;
wire [1:0] PT_F1L5_Plus_start;
wire [1:0] ME_F1F2_F3D5PHI3X1_start;
wire [1:0] TC_F1D5F2D5_proj_start;
wire [1:0] TE_F3D5PHI4X2_F4D5PHI3X2_start;
wire [1:0] VMS_F4D5PHI2X2n3_start;
wire [1:0] CM_F1F2_F4D5PHI1X1_start;
wire [1:0] ME_F3F4_F5D5PHI3X2_start;
wire [1:0] SP_F3D5PHI1X1_F4D5PHI1X1_start;
wire [1:0] VMPROJ_F3F4_F5D5PHI4X1_start;
wire [1:0] TE_F1D5PHI3X2_F2D5PHI2X2_start;
wire [1:0] VMPROJ_F1F2_F5D5PHI1X2_start;
wire [1:0] VMS_F1D5PHI3X1n3_start;
wire [1:0] ME_F1F2_F5D5PHI1X2_start;
wire [1:0] VMS_F2D5PHI2X1n2_start;
wire [1:0] ME_F3F4_F5D5PHI1X1_start;
wire [1:0] VMPROJ_F3F4_F5D5PHI3X1_start;
wire [1:0] VMPROJ_F1F2_F3D5PHI2X1_start;
wire [1:0] SD1_F4D5_start;
wire [1:0] TF_F1F2_start;
wire [1:0] ME_F3F4_F5D5PHI2X1_start;
wire [1:0] VMPROJ_F3F4_F1D5PHI4X2_start;
wire [1:0] TPROJ_ToMinus_F3D5F4D5_F2_start;
wire [1:0] VMS_F3D5PHI2X1n3_start;
wire [1:0] TE_F3D5PHI2X2_F4D5PHI2X2_start;
wire [1:0] TE_F3D5PHI3X2_F4D5PHI2X2_start;
wire [1:0] VMS_F3D5PHI3X1n4_start;
wire [1:0] MC_F3F4_F1D5_start;
wire [1:0] DR2_D5_start;
wire [1:0] PRD_F4D5_F1F2_start;
wire [1:0] ME_F1F2_F3D5PHI2X2_start;
wire [1:0] VMPROJ_F3F4_F1D5PHI1X2_start;
wire [1:0] FM_F1F2_F5_FromPlus_start;
wire [1:0] CM_F1F2_F5D5PHI1X1_start;
wire [1:0] VMS_F2D5PHI3X2n3_start;
wire [1:0] VMPROJ_F3F4_F1D5PHI3X2_start;
wire [1:0] VMPROJ_F3F4_F2D5PHI3X2_start;
wire [1:0] VMPROJ_F1F2_F4D5PHI2X2_start;
wire [1:0] VMPROJ_F1F2_F4D5PHI1X1_start;
wire [1:0] ME_F1F2_F5D5PHI2X2_start;
wire [1:0] VMS_F3D5PHI3X1n2_start;
wire [1:0] VMPROJ_F3F4_F2D5PHI1X1_start;
wire [1:0] TE_F1D5PHI4X2_F2D5PHI3X2_start;
wire [1:0] TPROJ_FromPlus_F4D5_F1F2_start;
wire [1:0] VMPROJ_F1F2_F4D5PHI3X1_start;
wire [1:0] TC_F3D5F4D5_proj_start;
wire [1:0] TE_F1D5PHI1X2_F2D5PHI1X2_start;
wire [1:0] FM_F1F2_F3D5_ToPlus_start;
wire [1:0] VMPROJ_F1F2_F3D5PHI4X1_start;
wire [1:0] ME_F3F4_F2D5PHI3X2_start;
wire [1:0] VMPROJ_F1F2_F5D5PHI4X1_start;
wire [1:0] VMS_F4D5PHI3X2n3_start;
wire [1:0] ME_F3F4_F1D5PHI2X1_start;
wire [1:0] VMS_F1D5PHI1X1n2_start;
wire [1:0] VMPROJ_F3F4_F1D5PHI2X1_start;
wire [1:0] SP_F1D5PHI1X1_F2D5PHI1X1_start;
wire [1:0] MT_FDSK_Plus_start;
wire [1:0] MC_F3F4_F2D5_start;
wire [1:0] ME_F1F2_F4D5PHI1X2_start;
wire [1:0] TE_F3D5PHI4X1_F4D5PHI3X1_start;
wire [1:0] ME_F3F4_F2D5PHI1X2_start;
wire [1:0] TE_F1D5PHI3X1_F2D5PHI2X1_start;
wire [1:0] ME_F1F2_F4D5PHI3X2_start;
wire [1:0] VMPROJ_F3F4_F5D5PHI2X2_start;
wire [1:0] VMS_F1D5PHI1X1n1_start;
wire [1:0] VMPROJ_F3F4_F5D5PHI1X2_start;
wire [1:0] VMPROJ_F3F4_F1D5PHI3X1_start;
wire [1:0] VMPROJ_F1F2_F5D5PHI1X1_start;
wire [1:0] VMS_F1D5PHI4X1n2_start;
wire [1:0] ME_F3F4_F5D5PHI4X2_start;
wire [1:0] VMS_F2D5PHI1X2n4_start;
wire [1:0] TPROJ_FromPlus_F5D5_F1F2_start;
wire [1:0] MT_FDSK_Minus_start;
wire [1:0] VMPROJ_F3F4_F1D5PHI1X1_start;
wire [1:0] VMS_F2D5PHI1X2n3_start;
wire [1:0] ME_F1F2_F5D5PHI1X1_start;
wire [1:0] VMS_F2D5PHI1X1n2_start;
wire [1:0] PT_L2L4F2_Plus_start;
wire [1:0] PRD_F2D5_F3F4_start;
wire [1:0] ME_F1F2_F3D5PHI1X1_start;
wire [1:0] TPROJ_ToMinus_F3D5F4D5_F1_start;
wire [1:0] PT_L2L4F2_Minus_start;
wire [1:0] PRD_F3D5_F1F2_start;
wire [1:0] MC_F1F2_F5D5_start;
wire [1:0] TE_F3D5PHI2X1_F4D5PHI1X2_start;
wire [1:0] VMS_F3D5PHI2X1n4_start;
wire [1:0] VMPROJ_F3F4_F2D5PHI1X2_start;
wire [1:0] ME_F1F2_F5D5PHI4X1_start;
wire [1:0] TE_F1D5PHI3X1_F2D5PHI3X1_start;
wire [1:0] ME_F3F4_F2D5PHI1X1_start;
wire [1:0] MC_F3F4_F5D5_start;
wire [1:0] VMPROJ_F3F4_F5D5PHI2X1_start;
wire [1:0] DR1_D5_start;
wire [1:0] VMS_F1D5PHI3X1n2_start;
wire [1:0] VMPROJ_F3F4_F2D5PHI3X1_start;
wire [1:0] ME_F3F4_F5D5PHI2X2_start;
wire [1:0] VMPROJ_F3F4_F1D5PHI4X1_start;
wire [1:0] TE_F1D5PHI3X1_F2D5PHI3X2_start;
wire [1:0] VMPROJ_F3F4_F1D5PHI2X2_start;
wire [1:0] TE_F1D5PHI2X2_F2D5PHI1X2_start;
wire [1:0] TPROJ_ToMinus_F1D5F2D5_F5_start;
wire [1:0] ME_F3F4_F1D5PHI3X2_start;
wire [1:0] ME_F1F2_F3D5PHI4X2_start;
wire [1:0] TPROJ_ToPlus_F3D5F4D5_F2_start;
wire [1:0] VMS_F1D5PHI2X1n4_start;
wire [1:0] VMRD_F4D5_start;
wire [1:0] VMRD_F3D5_start;
wire [1:0] MC_F1F2_F3D5_start;
wire [1:0] FT_F3F4_start;
wire [1:0] VMPROJ_F1F2_F3D5PHI1X2_start;
wire [1:0] VMS_F2D5PHI2X2n3_start;
wire [1:0] TE_F1D5PHI4X1_F2D5PHI3X1_start;
wire [1:0] TE_F1D5PHI2X1_F2D5PHI1X1_start;
wire [1:0] TE_F3D5PHI3X1_F4D5PHI2X1_start;
wire [1:0] TC_F3D5F4D5_start;
wire [1:0] SD1_F1D5_start;
wire [1:0] ME_F1F2_F4D5PHI1X1_start;
wire [1:0] CM_F3F4_F2D5PHI1X1_start;
wire [1:0] PT_F1L5_Minus_start;
wire [1:0] VMPROJ_F3F4_F2D5PHI2X2_start;
wire [1:0] TE_F1D5PHI3X2_F2D5PHI3X2_start;
wire [1:0] VMS_F4D5PHI1X2n3_start;
wire [1:0] ME_F3F4_F2D5PHI2X2_start;
wire [1:0] PRD_F5D5_F1F2_start;
wire [1:0] VMS_F3D5PHI4X1n2_start;
wire [1:0] TE_F3D5PHI1X1_F4D5PHI1X1_start;
wire [1:0] ME_F3F4_F1D5PHI3X1_start;
wire [1:0] FT_F1F2_start;
wire [1:0] VMS_F3D5PHI1X1n2_start;
wire [1:0] TE_F3D5PHI2X1_F4D5PHI2X1_start;
wire [1:0] TPROJ_ToPlus_F1D5F2D5_F5_start;
wire [1:0] VMS_F2D5PHI3X2n4_start;
wire [1:0] ME_F1F2_F4D5PHI2X1_start;
wire [1:0] TPROJ_FromPlus_F2D5_F3F4_start;
wire [1:0] VMPROJ_F1F2_F5D5PHI2X1_start;
wire [1:0] TE_F1D5PHI3X1_F2D5PHI2X2_start;
wire [1:0] SD1_F5D5_start;
wire [1:0] ME_F1F2_F3D5PHI4X1_start;
wire [1:0] VMS_F4D5PHI3X2n4_start;
wire [1:0] VMS_F4D5PHI1X1n2_start;
wire [1:0] VMPROJ_F3F4_F5D5PHI4X2_start;
wire [1:0] VMS_F4D5PHI2X1n2_start;
wire [1:0] VMRD_F5D5_start;
wire [1:0] VMS_F2D5PHI2X2n4_start;
wire [1:0] TC_F1D5F2D5_start;
wire [1:0] TPROJ_FromPlus_F5D5_F3F4_start;
wire [1:0] VMS_F1D5PHI2X1n3_start;
wire [1:0] ME_F3F4_F5D5PHI4X1_start;
wire [1:0] VMS_F1D5PHI3X1n4_start;
wire [1:0] ME_F3F4_F5D5PHI1X2_start;
wire [1:0] TE_F3D5PHI3X1_F4D5PHI3X1_start;
wire [1:0] TE_F3D5PHI1X2_F4D5PHI1X2_start;
wire [1:0] ME_F1F2_F5D5PHI3X2_start;
wire [1:0] VMPROJ_F3F4_F5D5PHI3X2_start;
wire [1:0] VMPROJ_F1F2_F3D5PHI3X2_start;
wire [1:0] PRD_F5D5_F3F4_start;
wire [1:0] VMS_F4D5PHI2X2n4_start;
wire [1:0] ME_F3F4_F1D5PHI1X1_start;
wire [1:0] ME_F1F2_F3D5PHI3X2_start;
wire [1:0] TPROJ_FromPlus_F3D5_F1F2_start;
wire [1:0] TE_F1D5PHI2X1_F2D5PHI1X2_start;
wire [1:0] TE_F3D5PHI2X1_F4D5PHI2X2_start;
wire [1:0] PD_start;
wire [1:0] ME_F3F4_F1D5PHI4X2_start;
wire [1:0] TE_F1D5PHI2X1_F2D5PHI2X2_start;
wire [1:0] VMPROJ_F1F2_F4D5PHI2X1_start;
wire [1:0] TE_F3D5PHI2X1_F4D5PHI1X1_start;
wire [1:0] VMS_F1D5PHI2X1n2_start;
wire [1:0] TE_F3D5PHI3X1_F4D5PHI3X2_start;
wire [1:0] VMRD_F2D5_start;
wire [1:0] VMPROJ_F1F2_F5D5PHI2X2_start;
wire [1:0] ME_F3F4_F1D5PHI4X1_start;
wire [1:0] ME_F3F4_F1D5PHI2X2_start;
wire [1:0] ME_F3F4_F5D5PHI3X1_start;
wire [1:0] TE_F1D5PHI1X1_F2D5PHI1X2_start;
wire [1:0] VMS_F3D5PHI2X1n2_start;
wire [1:0] TE_F1D5PHI2X2_F2D5PHI2X2_start;
wire [1:0] ME_F1F2_F5D5PHI3X1_start;
wire [1:0] ME_F1F2_F4D5PHI2X2_start;
wire [1:0] TE_F3D5PHI3X2_F4D5PHI3X2_start;
wire [1:0] VMPROJ_F1F2_F5D5PHI4X2_start;
wire [1:0] VMPROJ_F1F2_F5D5PHI3X2_start;
wire [1:0] SD1_F2D5_start;
wire [1:0] VMPROJ_F1F2_F3D5PHI2X2_start;
wire [1:0] ME_F3F4_F2D5PHI3X1_start;
wire [1:0] FM_F1F2_F3D5_ToMinus_start;
wire [1:0] ME_F1F2_F3D5PHI1X2_start;
wire [1:0] VMPROJ_F3F4_F2D5PHI2X1_start;
wire [1:0] MC_F1F2_F4D5_start;
wire [1:0] VMS_F3D5PHI3X1n3_start;
wire [1:0] TPROJ_FromPlus_F1D5_F3F4_start;
wire [1:0] TPROJ_ToPlus_F1D5F2D5_F4_start;
wire [1:0] ME_F1F2_F5D5PHI4X2_start;
wire [1:0] TE_F1D5PHI2X1_F2D5PHI2X1_start;
wire [1:0] VMRD_F1D5_start;
wire [1:0] CM_F1F2_F3D5PHI1X1_start;
wire [1:0] TE_F3D5PHI3X1_F4D5PHI2X2_start;
wire [1:0] FM_F3F4_F5_FromPlus_start;
wire [1:0] CM_F3F4_F5D5PHI1X1_start;
wire [1:0] ME_F1F2_F4D5PHI3X1_start;
wire [1:0] VMPROJ_F1F2_F4D5PHI3X2_start;
wire [1:0] CM_F3F4_F1D5PHI1X1_start;
wire [1:0] ME_F3F4_F2D5PHI2X1_start;
wire [1:0] ME_F3F4_F1D5PHI1X2_start;
wire [1:0] PT_L1L6F4_Minus_start;
wire [1:0] PT_L3F3F5_Plus_start;
wire [1:0] TPROJ_ToMinus_F1D5F2D5_F4_start;
wire [1:0] VMS_F4D5PHI1X2n4_start;
wire [1:0] TE_F3D5PHI1X1_F4D5PHI1X2_start;
wire [1:0] TE_F3D5PHI4X1_F4D5PHI3X2_start;
wire [1:0] PT_L1L6F4_Plus_start;
wire [1:0] VMPROJ_F1F2_F3D5PHI4X2_start;
wire [1:0] VMS_F3D5PHI1X1n1_start;
wire [1:0] PRD_F1D5_F3F4_start;
wire [1:0] ME_F1F2_F3D5PHI2X1_start;
wire [1:0] TE_F1D5PHI1X1_F2D5PHI1X1_start;
wire [1:0] DR3_D5_start;
wire [1:0] ME_F1F2_F5D5PHI2X1_start;
wire [1:0] VMPROJ_F1F2_F3D5PHI1X1_start;
wire [1:0] VMS_F4D5PHI3X1n2_start;
wire [1:0] VMPROJ_F1F2_F3D5PHI3X1_start;
wire [1:0] VMPROJ_F3F4_F5D5PHI1X1_start;
wire [1:0] VMPROJ_F1F2_F4D5PHI1X2_start;
wire [1:0] TE_F3D5PHI2X2_F4D5PHI1X2_start;

wire [53:0] TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F5;
wire TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F5_wr_en;
wire [5:0] TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_F1D5F2D5_F5(
.data_in(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F5),
.enable(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F5_wr_en),
.number_out(TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_ToPlus_F1D5F2D5_F5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F5;
wire TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F5_wr_en;
wire [5:0] TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_F3D5F4D5_F5(
.data_in(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F5),
.enable(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F5_wr_en),
.number_out(TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_ToPlus_F3D5F4D5_F5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F3;
wire TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F3_wr_en;
wire [5:0] TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_F1D5F2D5_F3(
.data_in(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F3),
.enable(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F3_wr_en),
.number_out(TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_ToPlus_F1D5F2D5_F3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F2;
wire TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F2_wr_en;
wire [5:0] TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_F3D5F4D5_F2(
.data_in(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F2),
.enable(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F2_wr_en),
.number_out(TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_ToPlus_F3D5F4D5_F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F1;
wire TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F1_wr_en;
wire [5:0] TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus_number;
wire [9:0] TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_F3D5F4D5_F1(
.data_in(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F1),
.enable(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F1_wr_en),
.number_out(TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus_number),
.read_add(TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus_read_add),
.data_out(TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_ToPlus_F3D5F4D5_F1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F4;
wire TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F4_wr_en;
wire [5:0] TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_F1D5F2D5_F4(
.data_in(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F4),
.enable(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F4_wr_en),
.number_out(TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_ToPlus_F1D5F2D5_F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F5;
wire TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F5_wr_en;
wire [5:0] TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_F1D5F2D5_F5(
.data_in(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F5),
.enable(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F5_wr_en),
.number_out(TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_ToMinus_F1D5F2D5_F5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F5;
wire TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F5_wr_en;
wire [5:0] TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_F3D5F4D5_F5(
.data_in(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F5),
.enable(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F5_wr_en),
.number_out(TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_ToMinus_F3D5F4D5_F5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F3;
wire TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F3_wr_en;
wire [5:0] TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_F1D5F2D5_F3(
.data_in(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F3),
.enable(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F3_wr_en),
.number_out(TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_ToMinus_F1D5F2D5_F3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F2;
wire TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F2_wr_en;
wire [5:0] TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_F3D5F4D5_F2(
.data_in(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F2),
.enable(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F2_wr_en),
.number_out(TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_ToMinus_F3D5F4D5_F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F1;
wire TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F1_wr_en;
wire [5:0] TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus_number;
wire [9:0] TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_F3D5F4D5_F1(
.data_in(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F1),
.enable(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F1_wr_en),
.number_out(TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus_number),
.read_add(TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus_read_add),
.data_out(TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_ToMinus_F3D5F4D5_F1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F4;
wire TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F4_wr_en;
wire [5:0] TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_F1D5F2D5_F4(
.data_in(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F4),
.enable(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F4_wr_en),
.number_out(TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_ToMinus_F1D5F2D5_F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire IL1_D5_DR1_D5_read_en;
wire [35:0] IL1_D5_DR1_D5;
//wire IL1_D5_DR1_D5_empty;
InputLink  IL1_D5(
.data_in1(input_link1_reg1),
.data_in2(input_link1_reg2),
.read_en(IL1_D5_DR1_D5_read_en),
.data_out(IL1_D5_DR1_D5),
.empty(IL1_D5_DR1_D5_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire IL2_D5_DR2_D5_read_en;
wire [35:0] IL2_D5_DR2_D5;
//wire IL2_D5_DR2_D5_empty;
InputLink  IL2_D5(
.data_in1(input_link2_reg1),
.data_in2(input_link2_reg2),
.read_en(IL2_D5_DR2_D5_read_en),
.data_out(IL2_D5_DR2_D5),
.empty(IL2_D5_DR2_D5_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire IL3_D5_DR3_D5_read_en;
wire [35:0] IL3_D5_DR3_D5;
//wire IL3_D5_DR3_D5_empty;
InputLink  IL3_D5(
.data_in1(input_link3_reg1),
.data_in2(input_link3_reg2),
.read_en(IL3_D5_DR3_D5_read_en),
.data_out(IL3_D5_DR3_D5),
.empty(IL3_D5_DR3_D5_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR1_D5_SD1_F1D5;
wire DR1_D5_SD1_F1D5_wr_en;
wire [5:0] SD1_F1D5_VMRD_F1D5_number;
wire [8:0] SD1_F1D5_VMRD_F1D5_read_add;
wire [35:0] SD1_F1D5_VMRD_F1D5;
StubsByLayer  SD1_F1D5(
.data_in(DR1_D5_SD1_F1D5),
.enable(DR1_D5_SD1_F1D5_wr_en),
.number_out(SD1_F1D5_VMRD_F1D5_number),
.read_add(SD1_F1D5_VMRD_F1D5_read_add),
.data_out(SD1_F1D5_VMRD_F1D5),
.start(DR1_D5_start),
.done(SD1_F1D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR2_D5_SD2_F1D5;
wire DR2_D5_SD2_F1D5_wr_en;
wire [5:0] SD2_F1D5_VMRD_F1D5_number;
wire [8:0] SD2_F1D5_VMRD_F1D5_read_add;
wire [35:0] SD2_F1D5_VMRD_F1D5;
StubsByLayer  SD2_F1D5(
.data_in(DR2_D5_SD2_F1D5),
.enable(DR2_D5_SD2_F1D5_wr_en),
.number_out(SD2_F1D5_VMRD_F1D5_number),
.read_add(SD2_F1D5_VMRD_F1D5_read_add),
.data_out(SD2_F1D5_VMRD_F1D5),
.start(DR2_D5_start),
.done(SD2_F1D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR3_D5_SD3_F1D5;
wire DR3_D5_SD3_F1D5_wr_en;
wire [5:0] SD3_F1D5_VMRD_F1D5_number;
wire [8:0] SD3_F1D5_VMRD_F1D5_read_add;
wire [35:0] SD3_F1D5_VMRD_F1D5;
StubsByLayer  SD3_F1D5(
.data_in(DR3_D5_SD3_F1D5),
.enable(DR3_D5_SD3_F1D5_wr_en),
.number_out(SD3_F1D5_VMRD_F1D5_number),
.read_add(SD3_F1D5_VMRD_F1D5_read_add),
.data_out(SD3_F1D5_VMRD_F1D5),
.start(DR3_D5_start),
.done(SD3_F1D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR1_D5_SD1_F2D5;
wire DR1_D5_SD1_F2D5_wr_en;
wire [5:0] SD1_F2D5_VMRD_F2D5_number;
wire [8:0] SD1_F2D5_VMRD_F2D5_read_add;
wire [35:0] SD1_F2D5_VMRD_F2D5;
StubsByLayer  SD1_F2D5(
.data_in(DR1_D5_SD1_F2D5),
.enable(DR1_D5_SD1_F2D5_wr_en),
.number_out(SD1_F2D5_VMRD_F2D5_number),
.read_add(SD1_F2D5_VMRD_F2D5_read_add),
.data_out(SD1_F2D5_VMRD_F2D5),
.start(DR1_D5_start),
.done(SD1_F2D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR2_D5_SD2_F2D5;
wire DR2_D5_SD2_F2D5_wr_en;
wire [5:0] SD2_F2D5_VMRD_F2D5_number;
wire [8:0] SD2_F2D5_VMRD_F2D5_read_add;
wire [35:0] SD2_F2D5_VMRD_F2D5;
StubsByLayer  SD2_F2D5(
.data_in(DR2_D5_SD2_F2D5),
.enable(DR2_D5_SD2_F2D5_wr_en),
.number_out(SD2_F2D5_VMRD_F2D5_number),
.read_add(SD2_F2D5_VMRD_F2D5_read_add),
.data_out(SD2_F2D5_VMRD_F2D5),
.start(DR2_D5_start),
.done(SD2_F2D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR3_D5_SD3_F2D5;
wire DR3_D5_SD3_F2D5_wr_en;
wire [5:0] SD3_F2D5_VMRD_F2D5_number;
wire [8:0] SD3_F2D5_VMRD_F2D5_read_add;
wire [35:0] SD3_F2D5_VMRD_F2D5;
StubsByLayer  SD3_F2D5(
.data_in(DR3_D5_SD3_F2D5),
.enable(DR3_D5_SD3_F2D5_wr_en),
.number_out(SD3_F2D5_VMRD_F2D5_number),
.read_add(SD3_F2D5_VMRD_F2D5_read_add),
.data_out(SD3_F2D5_VMRD_F2D5),
.start(DR3_D5_start),
.done(SD3_F2D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR1_D5_SD1_F3D5;
wire DR1_D5_SD1_F3D5_wr_en;
wire [5:0] SD1_F3D5_VMRD_F3D5_number;
wire [8:0] SD1_F3D5_VMRD_F3D5_read_add;
wire [35:0] SD1_F3D5_VMRD_F3D5;
StubsByLayer  SD1_F3D5(
.data_in(DR1_D5_SD1_F3D5),
.enable(DR1_D5_SD1_F3D5_wr_en),
.number_out(SD1_F3D5_VMRD_F3D5_number),
.read_add(SD1_F3D5_VMRD_F3D5_read_add),
.data_out(SD1_F3D5_VMRD_F3D5),
.start(DR1_D5_start),
.done(SD1_F3D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR2_D5_SD2_F3D5;
wire DR2_D5_SD2_F3D5_wr_en;
wire [5:0] SD2_F3D5_VMRD_F3D5_number;
wire [8:0] SD2_F3D5_VMRD_F3D5_read_add;
wire [35:0] SD2_F3D5_VMRD_F3D5;
StubsByLayer  SD2_F3D5(
.data_in(DR2_D5_SD2_F3D5),
.enable(DR2_D5_SD2_F3D5_wr_en),
.number_out(SD2_F3D5_VMRD_F3D5_number),
.read_add(SD2_F3D5_VMRD_F3D5_read_add),
.data_out(SD2_F3D5_VMRD_F3D5),
.start(DR2_D5_start),
.done(SD2_F3D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR3_D5_SD3_F3D5;
wire DR3_D5_SD3_F3D5_wr_en;
wire [5:0] SD3_F3D5_VMRD_F3D5_number;
wire [8:0] SD3_F3D5_VMRD_F3D5_read_add;
wire [35:0] SD3_F3D5_VMRD_F3D5;
StubsByLayer  SD3_F3D5(
.data_in(DR3_D5_SD3_F3D5),
.enable(DR3_D5_SD3_F3D5_wr_en),
.number_out(SD3_F3D5_VMRD_F3D5_number),
.read_add(SD3_F3D5_VMRD_F3D5_read_add),
.data_out(SD3_F3D5_VMRD_F3D5),
.start(DR3_D5_start),
.done(SD3_F3D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR1_D5_SD1_F4D5;
wire DR1_D5_SD1_F4D5_wr_en;
wire [5:0] SD1_F4D5_VMRD_F4D5_number;
wire [8:0] SD1_F4D5_VMRD_F4D5_read_add;
wire [35:0] SD1_F4D5_VMRD_F4D5;
StubsByLayer  SD1_F4D5(
.data_in(DR1_D5_SD1_F4D5),
.enable(DR1_D5_SD1_F4D5_wr_en),
.number_out(SD1_F4D5_VMRD_F4D5_number),
.read_add(SD1_F4D5_VMRD_F4D5_read_add),
.data_out(SD1_F4D5_VMRD_F4D5),
.start(DR1_D5_start),
.done(SD1_F4D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR2_D5_SD2_F4D5;
wire DR2_D5_SD2_F4D5_wr_en;
wire [5:0] SD2_F4D5_VMRD_F4D5_number;
wire [8:0] SD2_F4D5_VMRD_F4D5_read_add;
wire [35:0] SD2_F4D5_VMRD_F4D5;
StubsByLayer  SD2_F4D5(
.data_in(DR2_D5_SD2_F4D5),
.enable(DR2_D5_SD2_F4D5_wr_en),
.number_out(SD2_F4D5_VMRD_F4D5_number),
.read_add(SD2_F4D5_VMRD_F4D5_read_add),
.data_out(SD2_F4D5_VMRD_F4D5),
.start(DR2_D5_start),
.done(SD2_F4D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR3_D5_SD3_F4D5;
wire DR3_D5_SD3_F4D5_wr_en;
wire [5:0] SD3_F4D5_VMRD_F4D5_number;
wire [8:0] SD3_F4D5_VMRD_F4D5_read_add;
wire [35:0] SD3_F4D5_VMRD_F4D5;
StubsByLayer  SD3_F4D5(
.data_in(DR3_D5_SD3_F4D5),
.enable(DR3_D5_SD3_F4D5_wr_en),
.number_out(SD3_F4D5_VMRD_F4D5_number),
.read_add(SD3_F4D5_VMRD_F4D5_read_add),
.data_out(SD3_F4D5_VMRD_F4D5),
.start(DR3_D5_start),
.done(SD3_F4D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR1_D5_SD1_F5D5;
wire DR1_D5_SD1_F5D5_wr_en;
wire [5:0] SD1_F5D5_VMRD_F5D5_number;
wire [8:0] SD1_F5D5_VMRD_F5D5_read_add;
wire [35:0] SD1_F5D5_VMRD_F5D5;
StubsByLayer  SD1_F5D5(
.data_in(DR1_D5_SD1_F5D5),
.enable(DR1_D5_SD1_F5D5_wr_en),
.number_out(SD1_F5D5_VMRD_F5D5_number),
.read_add(SD1_F5D5_VMRD_F5D5_read_add),
.data_out(SD1_F5D5_VMRD_F5D5),
.start(DR1_D5_start),
.done(SD1_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR2_D5_SD2_F5D5;
wire DR2_D5_SD2_F5D5_wr_en;
wire [5:0] SD2_F5D5_VMRD_F5D5_number;
wire [8:0] SD2_F5D5_VMRD_F5D5_read_add;
wire [35:0] SD2_F5D5_VMRD_F5D5;
StubsByLayer  SD2_F5D5(
.data_in(DR2_D5_SD2_F5D5),
.enable(DR2_D5_SD2_F5D5_wr_en),
.number_out(SD2_F5D5_VMRD_F5D5_number),
.read_add(SD2_F5D5_VMRD_F5D5_read_add),
.data_out(SD2_F5D5_VMRD_F5D5),
.start(DR2_D5_start),
.done(SD2_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] DR3_D5_SD3_F5D5;
wire DR3_D5_SD3_F5D5_wr_en;
wire [5:0] SD3_F5D5_VMRD_F5D5_number;
wire [8:0] SD3_F5D5_VMRD_F5D5_read_add;
wire [35:0] SD3_F5D5_VMRD_F5D5;
StubsByLayer  SD3_F5D5(
.data_in(DR3_D5_SD3_F5D5),
.enable(DR3_D5_SD3_F5D5_wr_en),
.number_out(SD3_F5D5_VMRD_F5D5_number),
.read_add(SD3_F5D5_VMRD_F5D5_read_add),
.data_out(SD3_F5D5_VMRD_F5D5),
.start(DR3_D5_start),
.done(SD3_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI1X1n1;
wire VMRD_F1D5_VMS_F1D5PHI1X1n1_wr_en;
wire [5:0] VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_number;
wire [10:0] VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_read_add;
wire [18:0] VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1;
VMStubs #("Tracklet") VMS_F1D5PHI1X1n1(
.data_in(VMRD_F1D5_VMS_F1D5PHI1X1n1),
.enable(VMRD_F1D5_VMS_F1D5PHI1X1n1_wr_en),
.number_out(VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_number),
.read_add(VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_read_add),
.data_out(VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI1X1n1;
wire VMRD_F2D5_VMS_F2D5PHI1X1n1_wr_en;
wire [5:0] VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_number;
wire [10:0] VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_read_add;
wire [18:0] VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1;
VMStubs #("Tracklet") VMS_F2D5PHI1X1n1(
.data_in(VMRD_F2D5_VMS_F2D5PHI1X1n1),
.enable(VMRD_F2D5_VMS_F2D5PHI1X1n1_wr_en),
.number_out(VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_number),
.read_add(VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_read_add),
.data_out(VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI2X1n1;
wire VMRD_F1D5_VMS_F1D5PHI2X1n1_wr_en;
wire [5:0] VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1_number;
wire [10:0] VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1_read_add;
wire [18:0] VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1;
VMStubs #("Tracklet") VMS_F1D5PHI2X1n1(
.data_in(VMRD_F1D5_VMS_F1D5PHI2X1n1),
.enable(VMRD_F1D5_VMS_F1D5PHI2X1n1_wr_en),
.number_out(VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1_number),
.read_add(VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1_read_add),
.data_out(VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI1X1n2;
wire VMRD_F2D5_VMS_F2D5PHI1X1n2_wr_en;
wire [5:0] VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1_number;
wire [10:0] VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1_read_add;
wire [18:0] VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1;
VMStubs #("Tracklet") VMS_F2D5PHI1X1n2(
.data_in(VMRD_F2D5_VMS_F2D5PHI1X1n2),
.enable(VMRD_F2D5_VMS_F2D5PHI1X1n2_wr_en),
.number_out(VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1_number),
.read_add(VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1_read_add),
.data_out(VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI2X1n2;
wire VMRD_F1D5_VMS_F1D5PHI2X1n2_wr_en;
wire [5:0] VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1_number;
wire [10:0] VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1_read_add;
wire [18:0] VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1;
VMStubs #("Tracklet") VMS_F1D5PHI2X1n2(
.data_in(VMRD_F1D5_VMS_F1D5PHI2X1n2),
.enable(VMRD_F1D5_VMS_F1D5PHI2X1n2_wr_en),
.number_out(VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1_number),
.read_add(VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1_read_add),
.data_out(VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI2X1n1;
wire VMRD_F2D5_VMS_F2D5PHI2X1n1_wr_en;
wire [5:0] VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1_number;
wire [10:0] VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1_read_add;
wire [18:0] VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1;
VMStubs #("Tracklet") VMS_F2D5PHI2X1n1(
.data_in(VMRD_F2D5_VMS_F2D5PHI2X1n1),
.enable(VMRD_F2D5_VMS_F2D5PHI2X1n1_wr_en),
.number_out(VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1_number),
.read_add(VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1_read_add),
.data_out(VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI3X1n1;
wire VMRD_F1D5_VMS_F1D5PHI3X1n1_wr_en;
wire [5:0] VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1_number;
wire [10:0] VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1_read_add;
wire [18:0] VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1;
VMStubs #("Tracklet") VMS_F1D5PHI3X1n1(
.data_in(VMRD_F1D5_VMS_F1D5PHI3X1n1),
.enable(VMRD_F1D5_VMS_F1D5PHI3X1n1_wr_en),
.number_out(VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1_number),
.read_add(VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1_read_add),
.data_out(VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI2X1n2;
wire VMRD_F2D5_VMS_F2D5PHI2X1n2_wr_en;
wire [5:0] VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1_number;
wire [10:0] VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1_read_add;
wire [18:0] VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1;
VMStubs #("Tracklet") VMS_F2D5PHI2X1n2(
.data_in(VMRD_F2D5_VMS_F2D5PHI2X1n2),
.enable(VMRD_F2D5_VMS_F2D5PHI2X1n2_wr_en),
.number_out(VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1_number),
.read_add(VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1_read_add),
.data_out(VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI3X1n2;
wire VMRD_F1D5_VMS_F1D5PHI3X1n2_wr_en;
wire [5:0] VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1_number;
wire [10:0] VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1_read_add;
wire [18:0] VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1;
VMStubs #("Tracklet") VMS_F1D5PHI3X1n2(
.data_in(VMRD_F1D5_VMS_F1D5PHI3X1n2),
.enable(VMRD_F1D5_VMS_F1D5PHI3X1n2_wr_en),
.number_out(VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1_number),
.read_add(VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1_read_add),
.data_out(VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI3X1n1;
wire VMRD_F2D5_VMS_F2D5PHI3X1n1_wr_en;
wire [5:0] VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1_number;
wire [10:0] VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1_read_add;
wire [18:0] VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1;
VMStubs #("Tracklet") VMS_F2D5PHI3X1n1(
.data_in(VMRD_F2D5_VMS_F2D5PHI3X1n1),
.enable(VMRD_F2D5_VMS_F2D5PHI3X1n1_wr_en),
.number_out(VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1_number),
.read_add(VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1_read_add),
.data_out(VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI4X1n1;
wire VMRD_F1D5_VMS_F1D5PHI4X1n1_wr_en;
wire [5:0] VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1_number;
wire [10:0] VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1_read_add;
wire [18:0] VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1;
VMStubs #("Tracklet") VMS_F1D5PHI4X1n1(
.data_in(VMRD_F1D5_VMS_F1D5PHI4X1n1),
.enable(VMRD_F1D5_VMS_F1D5PHI4X1n1_wr_en),
.number_out(VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1_number),
.read_add(VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1_read_add),
.data_out(VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI3X1n2;
wire VMRD_F2D5_VMS_F2D5PHI3X1n2_wr_en;
wire [5:0] VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1_number;
wire [10:0] VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1_read_add;
wire [18:0] VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1;
VMStubs #("Tracklet") VMS_F2D5PHI3X1n2(
.data_in(VMRD_F2D5_VMS_F2D5PHI3X1n2),
.enable(VMRD_F2D5_VMS_F2D5PHI3X1n2_wr_en),
.number_out(VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1_number),
.read_add(VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1_read_add),
.data_out(VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI1X1n2;
wire VMRD_F1D5_VMS_F1D5PHI1X1n2_wr_en;
wire [5:0] VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2_number;
wire [10:0] VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2_read_add;
wire [18:0] VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2;
VMStubs #("Tracklet") VMS_F1D5PHI1X1n2(
.data_in(VMRD_F1D5_VMS_F1D5PHI1X1n2),
.enable(VMRD_F1D5_VMS_F1D5PHI1X1n2_wr_en),
.number_out(VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2_number),
.read_add(VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2_read_add),
.data_out(VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI1X2n1;
wire VMRD_F2D5_VMS_F2D5PHI1X2n1_wr_en;
wire [5:0] VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2_number;
wire [10:0] VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2_read_add;
wire [18:0] VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2;
VMStubs #("Tracklet") VMS_F2D5PHI1X2n1(
.data_in(VMRD_F2D5_VMS_F2D5PHI1X2n1),
.enable(VMRD_F2D5_VMS_F2D5PHI1X2n1_wr_en),
.number_out(VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2_number),
.read_add(VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2_read_add),
.data_out(VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI2X1n3;
wire VMRD_F1D5_VMS_F1D5PHI2X1n3_wr_en;
wire [5:0] VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2_number;
wire [10:0] VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2_read_add;
wire [18:0] VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2;
VMStubs #("Tracklet") VMS_F1D5PHI2X1n3(
.data_in(VMRD_F1D5_VMS_F1D5PHI2X1n3),
.enable(VMRD_F1D5_VMS_F1D5PHI2X1n3_wr_en),
.number_out(VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2_number),
.read_add(VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2_read_add),
.data_out(VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI1X2n2;
wire VMRD_F2D5_VMS_F2D5PHI1X2n2_wr_en;
wire [5:0] VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2_number;
wire [10:0] VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2_read_add;
wire [18:0] VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2;
VMStubs #("Tracklet") VMS_F2D5PHI1X2n2(
.data_in(VMRD_F2D5_VMS_F2D5PHI1X2n2),
.enable(VMRD_F2D5_VMS_F2D5PHI1X2n2_wr_en),
.number_out(VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2_number),
.read_add(VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2_read_add),
.data_out(VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI2X1n4;
wire VMRD_F1D5_VMS_F1D5PHI2X1n4_wr_en;
wire [5:0] VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2_number;
wire [10:0] VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2_read_add;
wire [18:0] VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2;
VMStubs #("Tracklet") VMS_F1D5PHI2X1n4(
.data_in(VMRD_F1D5_VMS_F1D5PHI2X1n4),
.enable(VMRD_F1D5_VMS_F1D5PHI2X1n4_wr_en),
.number_out(VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2_number),
.read_add(VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2_read_add),
.data_out(VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI2X2n1;
wire VMRD_F2D5_VMS_F2D5PHI2X2n1_wr_en;
wire [5:0] VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2_number;
wire [10:0] VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2_read_add;
wire [18:0] VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2;
VMStubs #("Tracklet") VMS_F2D5PHI2X2n1(
.data_in(VMRD_F2D5_VMS_F2D5PHI2X2n1),
.enable(VMRD_F2D5_VMS_F2D5PHI2X2n1_wr_en),
.number_out(VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2_number),
.read_add(VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2_read_add),
.data_out(VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI3X1n3;
wire VMRD_F1D5_VMS_F1D5PHI3X1n3_wr_en;
wire [5:0] VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2_number;
wire [10:0] VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2_read_add;
wire [18:0] VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2;
VMStubs #("Tracklet") VMS_F1D5PHI3X1n3(
.data_in(VMRD_F1D5_VMS_F1D5PHI3X1n3),
.enable(VMRD_F1D5_VMS_F1D5PHI3X1n3_wr_en),
.number_out(VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2_number),
.read_add(VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2_read_add),
.data_out(VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI2X2n2;
wire VMRD_F2D5_VMS_F2D5PHI2X2n2_wr_en;
wire [5:0] VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2_number;
wire [10:0] VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2_read_add;
wire [18:0] VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2;
VMStubs #("Tracklet") VMS_F2D5PHI2X2n2(
.data_in(VMRD_F2D5_VMS_F2D5PHI2X2n2),
.enable(VMRD_F2D5_VMS_F2D5PHI2X2n2_wr_en),
.number_out(VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2_number),
.read_add(VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2_read_add),
.data_out(VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI3X1n4;
wire VMRD_F1D5_VMS_F1D5PHI3X1n4_wr_en;
wire [5:0] VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2_number;
wire [10:0] VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2_read_add;
wire [18:0] VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2;
VMStubs #("Tracklet") VMS_F1D5PHI3X1n4(
.data_in(VMRD_F1D5_VMS_F1D5PHI3X1n4),
.enable(VMRD_F1D5_VMS_F1D5PHI3X1n4_wr_en),
.number_out(VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2_number),
.read_add(VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2_read_add),
.data_out(VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI3X2n1;
wire VMRD_F2D5_VMS_F2D5PHI3X2n1_wr_en;
wire [5:0] VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2_number;
wire [10:0] VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2_read_add;
wire [18:0] VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2;
VMStubs #("Tracklet") VMS_F2D5PHI3X2n1(
.data_in(VMRD_F2D5_VMS_F2D5PHI3X2n1),
.enable(VMRD_F2D5_VMS_F2D5PHI3X2n1_wr_en),
.number_out(VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2_number),
.read_add(VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2_read_add),
.data_out(VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI4X1n2;
wire VMRD_F1D5_VMS_F1D5PHI4X1n2_wr_en;
wire [5:0] VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2_number;
wire [10:0] VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2_read_add;
wire [18:0] VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2;
VMStubs #("Tracklet") VMS_F1D5PHI4X1n2(
.data_in(VMRD_F1D5_VMS_F1D5PHI4X1n2),
.enable(VMRD_F1D5_VMS_F1D5PHI4X1n2_wr_en),
.number_out(VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2_number),
.read_add(VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2_read_add),
.data_out(VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI3X2n2;
wire VMRD_F2D5_VMS_F2D5PHI3X2n2_wr_en;
wire [5:0] VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2_number;
wire [10:0] VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2_read_add;
wire [18:0] VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2;
VMStubs #("Tracklet") VMS_F2D5PHI3X2n2(
.data_in(VMRD_F2D5_VMS_F2D5PHI3X2n2),
.enable(VMRD_F2D5_VMS_F2D5PHI3X2n2_wr_en),
.number_out(VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2_number),
.read_add(VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2_read_add),
.data_out(VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI1X2n1;
wire VMRD_F1D5_VMS_F1D5PHI1X2n1_wr_en;
wire [5:0] VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2_number;
wire [10:0] VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2_read_add;
wire [18:0] VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2;
VMStubs #("Tracklet") VMS_F1D5PHI1X2n1(
.data_in(VMRD_F1D5_VMS_F1D5PHI1X2n1),
.enable(VMRD_F1D5_VMS_F1D5PHI1X2n1_wr_en),
.number_out(VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2_number),
.read_add(VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2_read_add),
.data_out(VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI1X2n3;
wire VMRD_F2D5_VMS_F2D5PHI1X2n3_wr_en;
wire [5:0] VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2_number;
wire [10:0] VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2_read_add;
wire [18:0] VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2;
VMStubs #("Tracklet") VMS_F2D5PHI1X2n3(
.data_in(VMRD_F2D5_VMS_F2D5PHI1X2n3),
.enable(VMRD_F2D5_VMS_F2D5PHI1X2n3_wr_en),
.number_out(VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2_number),
.read_add(VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2_read_add),
.data_out(VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI2X2n1;
wire VMRD_F1D5_VMS_F1D5PHI2X2n1_wr_en;
wire [5:0] VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2_number;
wire [10:0] VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2_read_add;
wire [18:0] VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2;
VMStubs #("Tracklet") VMS_F1D5PHI2X2n1(
.data_in(VMRD_F1D5_VMS_F1D5PHI2X2n1),
.enable(VMRD_F1D5_VMS_F1D5PHI2X2n1_wr_en),
.number_out(VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2_number),
.read_add(VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2_read_add),
.data_out(VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI1X2n4;
wire VMRD_F2D5_VMS_F2D5PHI1X2n4_wr_en;
wire [5:0] VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2_number;
wire [10:0] VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2_read_add;
wire [18:0] VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2;
VMStubs #("Tracklet") VMS_F2D5PHI1X2n4(
.data_in(VMRD_F2D5_VMS_F2D5PHI1X2n4),
.enable(VMRD_F2D5_VMS_F2D5PHI1X2n4_wr_en),
.number_out(VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2_number),
.read_add(VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2_read_add),
.data_out(VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI2X2n2;
wire VMRD_F1D5_VMS_F1D5PHI2X2n2_wr_en;
wire [5:0] VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2_number;
wire [10:0] VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2_read_add;
wire [18:0] VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2;
VMStubs #("Tracklet") VMS_F1D5PHI2X2n2(
.data_in(VMRD_F1D5_VMS_F1D5PHI2X2n2),
.enable(VMRD_F1D5_VMS_F1D5PHI2X2n2_wr_en),
.number_out(VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2_number),
.read_add(VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2_read_add),
.data_out(VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI2X2n3;
wire VMRD_F2D5_VMS_F2D5PHI2X2n3_wr_en;
wire [5:0] VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2_number;
wire [10:0] VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2_read_add;
wire [18:0] VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2;
VMStubs #("Tracklet") VMS_F2D5PHI2X2n3(
.data_in(VMRD_F2D5_VMS_F2D5PHI2X2n3),
.enable(VMRD_F2D5_VMS_F2D5PHI2X2n3_wr_en),
.number_out(VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2_number),
.read_add(VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2_read_add),
.data_out(VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI3X2n1;
wire VMRD_F1D5_VMS_F1D5PHI3X2n1_wr_en;
wire [5:0] VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2_number;
wire [10:0] VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2_read_add;
wire [18:0] VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2;
VMStubs #("Tracklet") VMS_F1D5PHI3X2n1(
.data_in(VMRD_F1D5_VMS_F1D5PHI3X2n1),
.enable(VMRD_F1D5_VMS_F1D5PHI3X2n1_wr_en),
.number_out(VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2_number),
.read_add(VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2_read_add),
.data_out(VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI2X2n4;
wire VMRD_F2D5_VMS_F2D5PHI2X2n4_wr_en;
wire [5:0] VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2_number;
wire [10:0] VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2_read_add;
wire [18:0] VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2;
VMStubs #("Tracklet") VMS_F2D5PHI2X2n4(
.data_in(VMRD_F2D5_VMS_F2D5PHI2X2n4),
.enable(VMRD_F2D5_VMS_F2D5PHI2X2n4_wr_en),
.number_out(VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2_number),
.read_add(VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2_read_add),
.data_out(VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI3X2n2;
wire VMRD_F1D5_VMS_F1D5PHI3X2n2_wr_en;
wire [5:0] VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2_number;
wire [10:0] VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2_read_add;
wire [18:0] VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2;
VMStubs #("Tracklet") VMS_F1D5PHI3X2n2(
.data_in(VMRD_F1D5_VMS_F1D5PHI3X2n2),
.enable(VMRD_F1D5_VMS_F1D5PHI3X2n2_wr_en),
.number_out(VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2_number),
.read_add(VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2_read_add),
.data_out(VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI3X2n3;
wire VMRD_F2D5_VMS_F2D5PHI3X2n3_wr_en;
wire [5:0] VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2_number;
wire [10:0] VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2_read_add;
wire [18:0] VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2;
VMStubs #("Tracklet") VMS_F2D5PHI3X2n3(
.data_in(VMRD_F2D5_VMS_F2D5PHI3X2n3),
.enable(VMRD_F2D5_VMS_F2D5PHI3X2n3_wr_en),
.number_out(VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2_number),
.read_add(VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2_read_add),
.data_out(VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI4X2n1;
wire VMRD_F1D5_VMS_F1D5PHI4X2n1_wr_en;
wire [5:0] VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2_number;
wire [10:0] VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2_read_add;
wire [18:0] VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2;
VMStubs #("Tracklet") VMS_F1D5PHI4X2n1(
.data_in(VMRD_F1D5_VMS_F1D5PHI4X2n1),
.enable(VMRD_F1D5_VMS_F1D5PHI4X2n1_wr_en),
.number_out(VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2_number),
.read_add(VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2_read_add),
.data_out(VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI3X2n4;
wire VMRD_F2D5_VMS_F2D5PHI3X2n4_wr_en;
wire [5:0] VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2_number;
wire [10:0] VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2_read_add;
wire [18:0] VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2;
VMStubs #("Tracklet") VMS_F2D5PHI3X2n4(
.data_in(VMRD_F2D5_VMS_F2D5PHI3X2n4),
.enable(VMRD_F2D5_VMS_F2D5PHI3X2n4_wr_en),
.number_out(VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2_number),
.read_add(VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2_read_add),
.data_out(VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI1X1n1;
wire VMRD_F3D5_VMS_F3D5PHI1X1n1_wr_en;
wire [5:0] VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_number;
wire [10:0] VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_read_add;
wire [18:0] VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1;
VMStubs #("Tracklet") VMS_F3D5PHI1X1n1(
.data_in(VMRD_F3D5_VMS_F3D5PHI1X1n1),
.enable(VMRD_F3D5_VMS_F3D5PHI1X1n1_wr_en),
.number_out(VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_number),
.read_add(VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_read_add),
.data_out(VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI1X1n1;
wire VMRD_F4D5_VMS_F4D5PHI1X1n1_wr_en;
wire [5:0] VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_number;
wire [10:0] VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_read_add;
wire [18:0] VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1;
VMStubs #("Tracklet") VMS_F4D5PHI1X1n1(
.data_in(VMRD_F4D5_VMS_F4D5PHI1X1n1),
.enable(VMRD_F4D5_VMS_F4D5PHI1X1n1_wr_en),
.number_out(VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_number),
.read_add(VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_read_add),
.data_out(VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI2X1n1;
wire VMRD_F3D5_VMS_F3D5PHI2X1n1_wr_en;
wire [5:0] VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1_number;
wire [10:0] VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1_read_add;
wire [18:0] VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1;
VMStubs #("Tracklet") VMS_F3D5PHI2X1n1(
.data_in(VMRD_F3D5_VMS_F3D5PHI2X1n1),
.enable(VMRD_F3D5_VMS_F3D5PHI2X1n1_wr_en),
.number_out(VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1_number),
.read_add(VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1_read_add),
.data_out(VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI1X1n2;
wire VMRD_F4D5_VMS_F4D5PHI1X1n2_wr_en;
wire [5:0] VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1_number;
wire [10:0] VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1_read_add;
wire [18:0] VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1;
VMStubs #("Tracklet") VMS_F4D5PHI1X1n2(
.data_in(VMRD_F4D5_VMS_F4D5PHI1X1n2),
.enable(VMRD_F4D5_VMS_F4D5PHI1X1n2_wr_en),
.number_out(VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1_number),
.read_add(VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1_read_add),
.data_out(VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI2X1n2;
wire VMRD_F3D5_VMS_F3D5PHI2X1n2_wr_en;
wire [5:0] VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1_number;
wire [10:0] VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1_read_add;
wire [18:0] VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1;
VMStubs #("Tracklet") VMS_F3D5PHI2X1n2(
.data_in(VMRD_F3D5_VMS_F3D5PHI2X1n2),
.enable(VMRD_F3D5_VMS_F3D5PHI2X1n2_wr_en),
.number_out(VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1_number),
.read_add(VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1_read_add),
.data_out(VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI2X1n1;
wire VMRD_F4D5_VMS_F4D5PHI2X1n1_wr_en;
wire [5:0] VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1_number;
wire [10:0] VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1_read_add;
wire [18:0] VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1;
VMStubs #("Tracklet") VMS_F4D5PHI2X1n1(
.data_in(VMRD_F4D5_VMS_F4D5PHI2X1n1),
.enable(VMRD_F4D5_VMS_F4D5PHI2X1n1_wr_en),
.number_out(VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1_number),
.read_add(VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1_read_add),
.data_out(VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI3X1n1;
wire VMRD_F3D5_VMS_F3D5PHI3X1n1_wr_en;
wire [5:0] VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1_number;
wire [10:0] VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1_read_add;
wire [18:0] VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1;
VMStubs #("Tracklet") VMS_F3D5PHI3X1n1(
.data_in(VMRD_F3D5_VMS_F3D5PHI3X1n1),
.enable(VMRD_F3D5_VMS_F3D5PHI3X1n1_wr_en),
.number_out(VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1_number),
.read_add(VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1_read_add),
.data_out(VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI2X1n2;
wire VMRD_F4D5_VMS_F4D5PHI2X1n2_wr_en;
wire [5:0] VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1_number;
wire [10:0] VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1_read_add;
wire [18:0] VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1;
VMStubs #("Tracklet") VMS_F4D5PHI2X1n2(
.data_in(VMRD_F4D5_VMS_F4D5PHI2X1n2),
.enable(VMRD_F4D5_VMS_F4D5PHI2X1n2_wr_en),
.number_out(VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1_number),
.read_add(VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1_read_add),
.data_out(VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI3X1n2;
wire VMRD_F3D5_VMS_F3D5PHI3X1n2_wr_en;
wire [5:0] VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1_number;
wire [10:0] VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1_read_add;
wire [18:0] VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1;
VMStubs #("Tracklet") VMS_F3D5PHI3X1n2(
.data_in(VMRD_F3D5_VMS_F3D5PHI3X1n2),
.enable(VMRD_F3D5_VMS_F3D5PHI3X1n2_wr_en),
.number_out(VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1_number),
.read_add(VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1_read_add),
.data_out(VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI3X1n1;
wire VMRD_F4D5_VMS_F4D5PHI3X1n1_wr_en;
wire [5:0] VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1_number;
wire [10:0] VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1_read_add;
wire [18:0] VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1;
VMStubs #("Tracklet") VMS_F4D5PHI3X1n1(
.data_in(VMRD_F4D5_VMS_F4D5PHI3X1n1),
.enable(VMRD_F4D5_VMS_F4D5PHI3X1n1_wr_en),
.number_out(VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1_number),
.read_add(VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1_read_add),
.data_out(VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI4X1n1;
wire VMRD_F3D5_VMS_F3D5PHI4X1n1_wr_en;
wire [5:0] VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1_number;
wire [10:0] VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1_read_add;
wire [18:0] VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1;
VMStubs #("Tracklet") VMS_F3D5PHI4X1n1(
.data_in(VMRD_F3D5_VMS_F3D5PHI4X1n1),
.enable(VMRD_F3D5_VMS_F3D5PHI4X1n1_wr_en),
.number_out(VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1_number),
.read_add(VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1_read_add),
.data_out(VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI3X1n2;
wire VMRD_F4D5_VMS_F4D5PHI3X1n2_wr_en;
wire [5:0] VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1_number;
wire [10:0] VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1_read_add;
wire [18:0] VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1;
VMStubs #("Tracklet") VMS_F4D5PHI3X1n2(
.data_in(VMRD_F4D5_VMS_F4D5PHI3X1n2),
.enable(VMRD_F4D5_VMS_F4D5PHI3X1n2_wr_en),
.number_out(VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1_number),
.read_add(VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1_read_add),
.data_out(VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI1X1n2;
wire VMRD_F3D5_VMS_F3D5PHI1X1n2_wr_en;
wire [5:0] VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2_number;
wire [10:0] VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2_read_add;
wire [18:0] VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2;
VMStubs #("Tracklet") VMS_F3D5PHI1X1n2(
.data_in(VMRD_F3D5_VMS_F3D5PHI1X1n2),
.enable(VMRD_F3D5_VMS_F3D5PHI1X1n2_wr_en),
.number_out(VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2_number),
.read_add(VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2_read_add),
.data_out(VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI1X2n1;
wire VMRD_F4D5_VMS_F4D5PHI1X2n1_wr_en;
wire [5:0] VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2_number;
wire [10:0] VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2_read_add;
wire [18:0] VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2;
VMStubs #("Tracklet") VMS_F4D5PHI1X2n1(
.data_in(VMRD_F4D5_VMS_F4D5PHI1X2n1),
.enable(VMRD_F4D5_VMS_F4D5PHI1X2n1_wr_en),
.number_out(VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2_number),
.read_add(VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2_read_add),
.data_out(VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI2X1n3;
wire VMRD_F3D5_VMS_F3D5PHI2X1n3_wr_en;
wire [5:0] VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2_number;
wire [10:0] VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2_read_add;
wire [18:0] VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2;
VMStubs #("Tracklet") VMS_F3D5PHI2X1n3(
.data_in(VMRD_F3D5_VMS_F3D5PHI2X1n3),
.enable(VMRD_F3D5_VMS_F3D5PHI2X1n3_wr_en),
.number_out(VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2_number),
.read_add(VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2_read_add),
.data_out(VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI1X2n2;
wire VMRD_F4D5_VMS_F4D5PHI1X2n2_wr_en;
wire [5:0] VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2_number;
wire [10:0] VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2_read_add;
wire [18:0] VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2;
VMStubs #("Tracklet") VMS_F4D5PHI1X2n2(
.data_in(VMRD_F4D5_VMS_F4D5PHI1X2n2),
.enable(VMRD_F4D5_VMS_F4D5PHI1X2n2_wr_en),
.number_out(VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2_number),
.read_add(VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2_read_add),
.data_out(VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI2X1n4;
wire VMRD_F3D5_VMS_F3D5PHI2X1n4_wr_en;
wire [5:0] VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2_number;
wire [10:0] VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2_read_add;
wire [18:0] VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2;
VMStubs #("Tracklet") VMS_F3D5PHI2X1n4(
.data_in(VMRD_F3D5_VMS_F3D5PHI2X1n4),
.enable(VMRD_F3D5_VMS_F3D5PHI2X1n4_wr_en),
.number_out(VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2_number),
.read_add(VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2_read_add),
.data_out(VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI2X2n1;
wire VMRD_F4D5_VMS_F4D5PHI2X2n1_wr_en;
wire [5:0] VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2_number;
wire [10:0] VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2_read_add;
wire [18:0] VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2;
VMStubs #("Tracklet") VMS_F4D5PHI2X2n1(
.data_in(VMRD_F4D5_VMS_F4D5PHI2X2n1),
.enable(VMRD_F4D5_VMS_F4D5PHI2X2n1_wr_en),
.number_out(VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2_number),
.read_add(VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2_read_add),
.data_out(VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI3X1n3;
wire VMRD_F3D5_VMS_F3D5PHI3X1n3_wr_en;
wire [5:0] VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2_number;
wire [10:0] VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2_read_add;
wire [18:0] VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2;
VMStubs #("Tracklet") VMS_F3D5PHI3X1n3(
.data_in(VMRD_F3D5_VMS_F3D5PHI3X1n3),
.enable(VMRD_F3D5_VMS_F3D5PHI3X1n3_wr_en),
.number_out(VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2_number),
.read_add(VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2_read_add),
.data_out(VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI2X2n2;
wire VMRD_F4D5_VMS_F4D5PHI2X2n2_wr_en;
wire [5:0] VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2_number;
wire [10:0] VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2_read_add;
wire [18:0] VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2;
VMStubs #("Tracklet") VMS_F4D5PHI2X2n2(
.data_in(VMRD_F4D5_VMS_F4D5PHI2X2n2),
.enable(VMRD_F4D5_VMS_F4D5PHI2X2n2_wr_en),
.number_out(VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2_number),
.read_add(VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2_read_add),
.data_out(VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI3X1n4;
wire VMRD_F3D5_VMS_F3D5PHI3X1n4_wr_en;
wire [5:0] VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2_number;
wire [10:0] VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2_read_add;
wire [18:0] VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2;
VMStubs #("Tracklet") VMS_F3D5PHI3X1n4(
.data_in(VMRD_F3D5_VMS_F3D5PHI3X1n4),
.enable(VMRD_F3D5_VMS_F3D5PHI3X1n4_wr_en),
.number_out(VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2_number),
.read_add(VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2_read_add),
.data_out(VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI3X2n1;
wire VMRD_F4D5_VMS_F4D5PHI3X2n1_wr_en;
wire [5:0] VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2_number;
wire [10:0] VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2_read_add;
wire [18:0] VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2;
VMStubs #("Tracklet") VMS_F4D5PHI3X2n1(
.data_in(VMRD_F4D5_VMS_F4D5PHI3X2n1),
.enable(VMRD_F4D5_VMS_F4D5PHI3X2n1_wr_en),
.number_out(VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2_number),
.read_add(VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2_read_add),
.data_out(VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI4X1n2;
wire VMRD_F3D5_VMS_F3D5PHI4X1n2_wr_en;
wire [5:0] VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2_number;
wire [10:0] VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2_read_add;
wire [18:0] VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2;
VMStubs #("Tracklet") VMS_F3D5PHI4X1n2(
.data_in(VMRD_F3D5_VMS_F3D5PHI4X1n2),
.enable(VMRD_F3D5_VMS_F3D5PHI4X1n2_wr_en),
.number_out(VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2_number),
.read_add(VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2_read_add),
.data_out(VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI3X2n2;
wire VMRD_F4D5_VMS_F4D5PHI3X2n2_wr_en;
wire [5:0] VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2_number;
wire [10:0] VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2_read_add;
wire [18:0] VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2;
VMStubs #("Tracklet") VMS_F4D5PHI3X2n2(
.data_in(VMRD_F4D5_VMS_F4D5PHI3X2n2),
.enable(VMRD_F4D5_VMS_F4D5PHI3X2n2_wr_en),
.number_out(VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2_number),
.read_add(VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2_read_add),
.data_out(VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI1X2n1;
wire VMRD_F3D5_VMS_F3D5PHI1X2n1_wr_en;
wire [5:0] VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2_number;
wire [10:0] VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2_read_add;
wire [18:0] VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2;
VMStubs #("Tracklet") VMS_F3D5PHI1X2n1(
.data_in(VMRD_F3D5_VMS_F3D5PHI1X2n1),
.enable(VMRD_F3D5_VMS_F3D5PHI1X2n1_wr_en),
.number_out(VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2_number),
.read_add(VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2_read_add),
.data_out(VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI1X2n3;
wire VMRD_F4D5_VMS_F4D5PHI1X2n3_wr_en;
wire [5:0] VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2_number;
wire [10:0] VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2_read_add;
wire [18:0] VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2;
VMStubs #("Tracklet") VMS_F4D5PHI1X2n3(
.data_in(VMRD_F4D5_VMS_F4D5PHI1X2n3),
.enable(VMRD_F4D5_VMS_F4D5PHI1X2n3_wr_en),
.number_out(VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2_number),
.read_add(VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2_read_add),
.data_out(VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI2X2n1;
wire VMRD_F3D5_VMS_F3D5PHI2X2n1_wr_en;
wire [5:0] VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2_number;
wire [10:0] VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2_read_add;
wire [18:0] VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2;
VMStubs #("Tracklet") VMS_F3D5PHI2X2n1(
.data_in(VMRD_F3D5_VMS_F3D5PHI2X2n1),
.enable(VMRD_F3D5_VMS_F3D5PHI2X2n1_wr_en),
.number_out(VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2_number),
.read_add(VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2_read_add),
.data_out(VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI1X2n4;
wire VMRD_F4D5_VMS_F4D5PHI1X2n4_wr_en;
wire [5:0] VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2_number;
wire [10:0] VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2_read_add;
wire [18:0] VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2;
VMStubs #("Tracklet") VMS_F4D5PHI1X2n4(
.data_in(VMRD_F4D5_VMS_F4D5PHI1X2n4),
.enable(VMRD_F4D5_VMS_F4D5PHI1X2n4_wr_en),
.number_out(VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2_number),
.read_add(VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2_read_add),
.data_out(VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI2X2n2;
wire VMRD_F3D5_VMS_F3D5PHI2X2n2_wr_en;
wire [5:0] VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2_number;
wire [10:0] VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2_read_add;
wire [18:0] VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2;
VMStubs #("Tracklet") VMS_F3D5PHI2X2n2(
.data_in(VMRD_F3D5_VMS_F3D5PHI2X2n2),
.enable(VMRD_F3D5_VMS_F3D5PHI2X2n2_wr_en),
.number_out(VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2_number),
.read_add(VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2_read_add),
.data_out(VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI2X2n3;
wire VMRD_F4D5_VMS_F4D5PHI2X2n3_wr_en;
wire [5:0] VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2_number;
wire [10:0] VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2_read_add;
wire [18:0] VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2;
VMStubs #("Tracklet") VMS_F4D5PHI2X2n3(
.data_in(VMRD_F4D5_VMS_F4D5PHI2X2n3),
.enable(VMRD_F4D5_VMS_F4D5PHI2X2n3_wr_en),
.number_out(VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2_number),
.read_add(VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2_read_add),
.data_out(VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI3X2n1;
wire VMRD_F3D5_VMS_F3D5PHI3X2n1_wr_en;
wire [5:0] VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2_number;
wire [10:0] VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2_read_add;
wire [18:0] VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2;
VMStubs #("Tracklet") VMS_F3D5PHI3X2n1(
.data_in(VMRD_F3D5_VMS_F3D5PHI3X2n1),
.enable(VMRD_F3D5_VMS_F3D5PHI3X2n1_wr_en),
.number_out(VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2_number),
.read_add(VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2_read_add),
.data_out(VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI2X2n4;
wire VMRD_F4D5_VMS_F4D5PHI2X2n4_wr_en;
wire [5:0] VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2_number;
wire [10:0] VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2_read_add;
wire [18:0] VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2;
VMStubs #("Tracklet") VMS_F4D5PHI2X2n4(
.data_in(VMRD_F4D5_VMS_F4D5PHI2X2n4),
.enable(VMRD_F4D5_VMS_F4D5PHI2X2n4_wr_en),
.number_out(VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2_number),
.read_add(VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2_read_add),
.data_out(VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI3X2n2;
wire VMRD_F3D5_VMS_F3D5PHI3X2n2_wr_en;
wire [5:0] VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2_number;
wire [10:0] VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2_read_add;
wire [18:0] VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2;
VMStubs #("Tracklet") VMS_F3D5PHI3X2n2(
.data_in(VMRD_F3D5_VMS_F3D5PHI3X2n2),
.enable(VMRD_F3D5_VMS_F3D5PHI3X2n2_wr_en),
.number_out(VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2_number),
.read_add(VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2_read_add),
.data_out(VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI3X2n3;
wire VMRD_F4D5_VMS_F4D5PHI3X2n3_wr_en;
wire [5:0] VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2_number;
wire [10:0] VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2_read_add;
wire [18:0] VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2;
VMStubs #("Tracklet") VMS_F4D5PHI3X2n3(
.data_in(VMRD_F4D5_VMS_F4D5PHI3X2n3),
.enable(VMRD_F4D5_VMS_F4D5PHI3X2n3_wr_en),
.number_out(VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2_number),
.read_add(VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2_read_add),
.data_out(VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI4X2n1;
wire VMRD_F3D5_VMS_F3D5PHI4X2n1_wr_en;
wire [5:0] VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2_number;
wire [10:0] VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2_read_add;
wire [18:0] VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2;
VMStubs #("Tracklet") VMS_F3D5PHI4X2n1(
.data_in(VMRD_F3D5_VMS_F3D5PHI4X2n1),
.enable(VMRD_F3D5_VMS_F3D5PHI4X2n1_wr_en),
.number_out(VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2_number),
.read_add(VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2_read_add),
.data_out(VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI3X2n4;
wire VMRD_F4D5_VMS_F4D5PHI3X2n4_wr_en;
wire [5:0] VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2_number;
wire [10:0] VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2_read_add;
wire [18:0] VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2;
VMStubs #("Tracklet") VMS_F4D5PHI3X2n4(
.data_in(VMRD_F4D5_VMS_F4D5PHI3X2n4),
.enable(VMRD_F4D5_VMS_F4D5PHI3X2n4_wr_en),
.number_out(VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2_number),
.read_add(VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2_read_add),
.data_out(VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI1X1_F2D5PHI1X1_SP_F1D5PHI1X1_F2D5PHI1X1;
wire TE_F1D5PHI1X1_F2D5PHI1X1_SP_F1D5PHI1X1_F2D5PHI1X1_wr_en;
wire [5:0] SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI1X1_F2D5PHI1X1(
.data_in(TE_F1D5PHI1X1_F2D5PHI1X1_SP_F1D5PHI1X1_F2D5PHI1X1),
.enable(TE_F1D5PHI1X1_F2D5PHI1X1_SP_F1D5PHI1X1_F2D5PHI1X1_wr_en),
.number_out(SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5),
.start(TE_F1D5PHI1X1_F2D5PHI1X1_start),
.done(SP_F1D5PHI1X1_F2D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI2X1_F2D5PHI1X1_SP_F1D5PHI2X1_F2D5PHI1X1;
wire TE_F1D5PHI2X1_F2D5PHI1X1_SP_F1D5PHI2X1_F2D5PHI1X1_wr_en;
wire [5:0] SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI2X1_F2D5PHI1X1(
.data_in(TE_F1D5PHI2X1_F2D5PHI1X1_SP_F1D5PHI2X1_F2D5PHI1X1),
.enable(TE_F1D5PHI2X1_F2D5PHI1X1_SP_F1D5PHI2X1_F2D5PHI1X1_wr_en),
.number_out(SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5),
.start(TE_F1D5PHI2X1_F2D5PHI1X1_start),
.done(SP_F1D5PHI2X1_F2D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI2X1_F2D5PHI2X1_SP_F1D5PHI2X1_F2D5PHI2X1;
wire TE_F1D5PHI2X1_F2D5PHI2X1_SP_F1D5PHI2X1_F2D5PHI2X1_wr_en;
wire [5:0] SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI2X1_F2D5PHI2X1(
.data_in(TE_F1D5PHI2X1_F2D5PHI2X1_SP_F1D5PHI2X1_F2D5PHI2X1),
.enable(TE_F1D5PHI2X1_F2D5PHI2X1_SP_F1D5PHI2X1_F2D5PHI2X1_wr_en),
.number_out(SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5),
.start(TE_F1D5PHI2X1_F2D5PHI2X1_start),
.done(SP_F1D5PHI2X1_F2D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI3X1_F2D5PHI2X1_SP_F1D5PHI3X1_F2D5PHI2X1;
wire TE_F1D5PHI3X1_F2D5PHI2X1_SP_F1D5PHI3X1_F2D5PHI2X1_wr_en;
wire [5:0] SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI3X1_F2D5PHI2X1(
.data_in(TE_F1D5PHI3X1_F2D5PHI2X1_SP_F1D5PHI3X1_F2D5PHI2X1),
.enable(TE_F1D5PHI3X1_F2D5PHI2X1_SP_F1D5PHI3X1_F2D5PHI2X1_wr_en),
.number_out(SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5),
.start(TE_F1D5PHI3X1_F2D5PHI2X1_start),
.done(SP_F1D5PHI3X1_F2D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI3X1_F2D5PHI3X1_SP_F1D5PHI3X1_F2D5PHI3X1;
wire TE_F1D5PHI3X1_F2D5PHI3X1_SP_F1D5PHI3X1_F2D5PHI3X1_wr_en;
wire [5:0] SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI3X1_F2D5PHI3X1(
.data_in(TE_F1D5PHI3X1_F2D5PHI3X1_SP_F1D5PHI3X1_F2D5PHI3X1),
.enable(TE_F1D5PHI3X1_F2D5PHI3X1_SP_F1D5PHI3X1_F2D5PHI3X1_wr_en),
.number_out(SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5),
.start(TE_F1D5PHI3X1_F2D5PHI3X1_start),
.done(SP_F1D5PHI3X1_F2D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI4X1_F2D5PHI3X1_SP_F1D5PHI4X1_F2D5PHI3X1;
wire TE_F1D5PHI4X1_F2D5PHI3X1_SP_F1D5PHI4X1_F2D5PHI3X1_wr_en;
wire [5:0] SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI4X1_F2D5PHI3X1(
.data_in(TE_F1D5PHI4X1_F2D5PHI3X1_SP_F1D5PHI4X1_F2D5PHI3X1),
.enable(TE_F1D5PHI4X1_F2D5PHI3X1_SP_F1D5PHI4X1_F2D5PHI3X1_wr_en),
.number_out(SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5),
.start(TE_F1D5PHI4X1_F2D5PHI3X1_start),
.done(SP_F1D5PHI4X1_F2D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI1X1_F2D5PHI1X2_SP_F1D5PHI1X1_F2D5PHI1X2;
wire TE_F1D5PHI1X1_F2D5PHI1X2_SP_F1D5PHI1X1_F2D5PHI1X2_wr_en;
wire [5:0] SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI1X1_F2D5PHI1X2(
.data_in(TE_F1D5PHI1X1_F2D5PHI1X2_SP_F1D5PHI1X1_F2D5PHI1X2),
.enable(TE_F1D5PHI1X1_F2D5PHI1X2_SP_F1D5PHI1X1_F2D5PHI1X2_wr_en),
.number_out(SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5),
.start(TE_F1D5PHI1X1_F2D5PHI1X2_start),
.done(SP_F1D5PHI1X1_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI2X1_F2D5PHI1X2_SP_F1D5PHI2X1_F2D5PHI1X2;
wire TE_F1D5PHI2X1_F2D5PHI1X2_SP_F1D5PHI2X1_F2D5PHI1X2_wr_en;
wire [5:0] SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI2X1_F2D5PHI1X2(
.data_in(TE_F1D5PHI2X1_F2D5PHI1X2_SP_F1D5PHI2X1_F2D5PHI1X2),
.enable(TE_F1D5PHI2X1_F2D5PHI1X2_SP_F1D5PHI2X1_F2D5PHI1X2_wr_en),
.number_out(SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5),
.start(TE_F1D5PHI2X1_F2D5PHI1X2_start),
.done(SP_F1D5PHI2X1_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI2X1_F2D5PHI2X2_SP_F1D5PHI2X1_F2D5PHI2X2;
wire TE_F1D5PHI2X1_F2D5PHI2X2_SP_F1D5PHI2X1_F2D5PHI2X2_wr_en;
wire [5:0] SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI2X1_F2D5PHI2X2(
.data_in(TE_F1D5PHI2X1_F2D5PHI2X2_SP_F1D5PHI2X1_F2D5PHI2X2),
.enable(TE_F1D5PHI2X1_F2D5PHI2X2_SP_F1D5PHI2X1_F2D5PHI2X2_wr_en),
.number_out(SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5),
.start(TE_F1D5PHI2X1_F2D5PHI2X2_start),
.done(SP_F1D5PHI2X1_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI3X1_F2D5PHI2X2_SP_F1D5PHI3X1_F2D5PHI2X2;
wire TE_F1D5PHI3X1_F2D5PHI2X2_SP_F1D5PHI3X1_F2D5PHI2X2_wr_en;
wire [5:0] SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI3X1_F2D5PHI2X2(
.data_in(TE_F1D5PHI3X1_F2D5PHI2X2_SP_F1D5PHI3X1_F2D5PHI2X2),
.enable(TE_F1D5PHI3X1_F2D5PHI2X2_SP_F1D5PHI3X1_F2D5PHI2X2_wr_en),
.number_out(SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5),
.start(TE_F1D5PHI3X1_F2D5PHI2X2_start),
.done(SP_F1D5PHI3X1_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI3X1_F2D5PHI3X2_SP_F1D5PHI3X1_F2D5PHI3X2;
wire TE_F1D5PHI3X1_F2D5PHI3X2_SP_F1D5PHI3X1_F2D5PHI3X2_wr_en;
wire [5:0] SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI3X1_F2D5PHI3X2(
.data_in(TE_F1D5PHI3X1_F2D5PHI3X2_SP_F1D5PHI3X1_F2D5PHI3X2),
.enable(TE_F1D5PHI3X1_F2D5PHI3X2_SP_F1D5PHI3X1_F2D5PHI3X2_wr_en),
.number_out(SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5),
.start(TE_F1D5PHI3X1_F2D5PHI3X2_start),
.done(SP_F1D5PHI3X1_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI4X1_F2D5PHI3X2_SP_F1D5PHI4X1_F2D5PHI3X2;
wire TE_F1D5PHI4X1_F2D5PHI3X2_SP_F1D5PHI4X1_F2D5PHI3X2_wr_en;
wire [5:0] SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI4X1_F2D5PHI3X2(
.data_in(TE_F1D5PHI4X1_F2D5PHI3X2_SP_F1D5PHI4X1_F2D5PHI3X2),
.enable(TE_F1D5PHI4X1_F2D5PHI3X2_SP_F1D5PHI4X1_F2D5PHI3X2_wr_en),
.number_out(SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5),
.start(TE_F1D5PHI4X1_F2D5PHI3X2_start),
.done(SP_F1D5PHI4X1_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI1X2_F2D5PHI1X2_SP_F1D5PHI1X2_F2D5PHI1X2;
wire TE_F1D5PHI1X2_F2D5PHI1X2_SP_F1D5PHI1X2_F2D5PHI1X2_wr_en;
wire [5:0] SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI1X2_F2D5PHI1X2(
.data_in(TE_F1D5PHI1X2_F2D5PHI1X2_SP_F1D5PHI1X2_F2D5PHI1X2),
.enable(TE_F1D5PHI1X2_F2D5PHI1X2_SP_F1D5PHI1X2_F2D5PHI1X2_wr_en),
.number_out(SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5),
.start(TE_F1D5PHI1X2_F2D5PHI1X2_start),
.done(SP_F1D5PHI1X2_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI2X2_F2D5PHI1X2_SP_F1D5PHI2X2_F2D5PHI1X2;
wire TE_F1D5PHI2X2_F2D5PHI1X2_SP_F1D5PHI2X2_F2D5PHI1X2_wr_en;
wire [5:0] SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI2X2_F2D5PHI1X2(
.data_in(TE_F1D5PHI2X2_F2D5PHI1X2_SP_F1D5PHI2X2_F2D5PHI1X2),
.enable(TE_F1D5PHI2X2_F2D5PHI1X2_SP_F1D5PHI2X2_F2D5PHI1X2_wr_en),
.number_out(SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5),
.start(TE_F1D5PHI2X2_F2D5PHI1X2_start),
.done(SP_F1D5PHI2X2_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI2X2_F2D5PHI2X2_SP_F1D5PHI2X2_F2D5PHI2X2;
wire TE_F1D5PHI2X2_F2D5PHI2X2_SP_F1D5PHI2X2_F2D5PHI2X2_wr_en;
wire [5:0] SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI2X2_F2D5PHI2X2(
.data_in(TE_F1D5PHI2X2_F2D5PHI2X2_SP_F1D5PHI2X2_F2D5PHI2X2),
.enable(TE_F1D5PHI2X2_F2D5PHI2X2_SP_F1D5PHI2X2_F2D5PHI2X2_wr_en),
.number_out(SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5),
.start(TE_F1D5PHI2X2_F2D5PHI2X2_start),
.done(SP_F1D5PHI2X2_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI3X2_F2D5PHI2X2_SP_F1D5PHI3X2_F2D5PHI2X2;
wire TE_F1D5PHI3X2_F2D5PHI2X2_SP_F1D5PHI3X2_F2D5PHI2X2_wr_en;
wire [5:0] SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI3X2_F2D5PHI2X2(
.data_in(TE_F1D5PHI3X2_F2D5PHI2X2_SP_F1D5PHI3X2_F2D5PHI2X2),
.enable(TE_F1D5PHI3X2_F2D5PHI2X2_SP_F1D5PHI3X2_F2D5PHI2X2_wr_en),
.number_out(SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5),
.start(TE_F1D5PHI3X2_F2D5PHI2X2_start),
.done(SP_F1D5PHI3X2_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI3X2_F2D5PHI3X2_SP_F1D5PHI3X2_F2D5PHI3X2;
wire TE_F1D5PHI3X2_F2D5PHI3X2_SP_F1D5PHI3X2_F2D5PHI3X2_wr_en;
wire [5:0] SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI3X2_F2D5PHI3X2(
.data_in(TE_F1D5PHI3X2_F2D5PHI3X2_SP_F1D5PHI3X2_F2D5PHI3X2),
.enable(TE_F1D5PHI3X2_F2D5PHI3X2_SP_F1D5PHI3X2_F2D5PHI3X2_wr_en),
.number_out(SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5),
.start(TE_F1D5PHI3X2_F2D5PHI3X2_start),
.done(SP_F1D5PHI3X2_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F1D5PHI4X2_F2D5PHI3X2_SP_F1D5PHI4X2_F2D5PHI3X2;
wire TE_F1D5PHI4X2_F2D5PHI3X2_SP_F1D5PHI4X2_F2D5PHI3X2_wr_en;
wire [5:0] SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5_number;
wire [8:0] SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5_read_add;
wire [11:0] SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5;
StubPairs  SP_F1D5PHI4X2_F2D5PHI3X2(
.data_in(TE_F1D5PHI4X2_F2D5PHI3X2_SP_F1D5PHI4X2_F2D5PHI3X2),
.enable(TE_F1D5PHI4X2_F2D5PHI3X2_SP_F1D5PHI4X2_F2D5PHI3X2_wr_en),
.number_out(SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5_number),
.read_add(SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5_read_add),
.data_out(SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5),
.start(TE_F1D5PHI4X2_F2D5PHI3X2_start),
.done(SP_F1D5PHI4X2_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F1D5_AS_F1D5n1;
wire VMRD_F1D5_AS_F1D5n1_wr_en;
wire [10:0] AS_F1D5n1_TC_F1D5F2D5_read_add;
wire [35:0] AS_F1D5n1_TC_F1D5F2D5;
AllStubs  AS_F1D5n1(
.data_in(VMRD_F1D5_AS_F1D5n1),
.enable(VMRD_F1D5_AS_F1D5n1_wr_en),
.read_add(AS_F1D5n1_TC_F1D5F2D5_read_add),
.data_out(AS_F1D5n1_TC_F1D5F2D5),
.start(VMRD_F1D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F2D5_AS_F2D5n1;
wire VMRD_F2D5_AS_F2D5n1_wr_en;
wire [10:0] AS_F2D5n1_TC_F1D5F2D5_read_add;
wire [35:0] AS_F2D5n1_TC_F1D5F2D5;
AllStubs  AS_F2D5n1(
.data_in(VMRD_F2D5_AS_F2D5n1),
.enable(VMRD_F2D5_AS_F2D5n1_wr_en),
.read_add(AS_F2D5n1_TC_F1D5F2D5_read_add),
.data_out(AS_F2D5n1_TC_F1D5F2D5),
.start(VMRD_F2D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI1X1_F4D5PHI1X1_SP_F3D5PHI1X1_F4D5PHI1X1;
wire TE_F3D5PHI1X1_F4D5PHI1X1_SP_F3D5PHI1X1_F4D5PHI1X1_wr_en;
wire [5:0] SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI1X1_F4D5PHI1X1(
.data_in(TE_F3D5PHI1X1_F4D5PHI1X1_SP_F3D5PHI1X1_F4D5PHI1X1),
.enable(TE_F3D5PHI1X1_F4D5PHI1X1_SP_F3D5PHI1X1_F4D5PHI1X1_wr_en),
.number_out(SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5),
.start(TE_F3D5PHI1X1_F4D5PHI1X1_start),
.done(SP_F3D5PHI1X1_F4D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI2X1_F4D5PHI1X1_SP_F3D5PHI2X1_F4D5PHI1X1;
wire TE_F3D5PHI2X1_F4D5PHI1X1_SP_F3D5PHI2X1_F4D5PHI1X1_wr_en;
wire [5:0] SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI2X1_F4D5PHI1X1(
.data_in(TE_F3D5PHI2X1_F4D5PHI1X1_SP_F3D5PHI2X1_F4D5PHI1X1),
.enable(TE_F3D5PHI2X1_F4D5PHI1X1_SP_F3D5PHI2X1_F4D5PHI1X1_wr_en),
.number_out(SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5),
.start(TE_F3D5PHI2X1_F4D5PHI1X1_start),
.done(SP_F3D5PHI2X1_F4D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI2X1_F4D5PHI2X1_SP_F3D5PHI2X1_F4D5PHI2X1;
wire TE_F3D5PHI2X1_F4D5PHI2X1_SP_F3D5PHI2X1_F4D5PHI2X1_wr_en;
wire [5:0] SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI2X1_F4D5PHI2X1(
.data_in(TE_F3D5PHI2X1_F4D5PHI2X1_SP_F3D5PHI2X1_F4D5PHI2X1),
.enable(TE_F3D5PHI2X1_F4D5PHI2X1_SP_F3D5PHI2X1_F4D5PHI2X1_wr_en),
.number_out(SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5),
.start(TE_F3D5PHI2X1_F4D5PHI2X1_start),
.done(SP_F3D5PHI2X1_F4D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI3X1_F4D5PHI2X1_SP_F3D5PHI3X1_F4D5PHI2X1;
wire TE_F3D5PHI3X1_F4D5PHI2X1_SP_F3D5PHI3X1_F4D5PHI2X1_wr_en;
wire [5:0] SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI3X1_F4D5PHI2X1(
.data_in(TE_F3D5PHI3X1_F4D5PHI2X1_SP_F3D5PHI3X1_F4D5PHI2X1),
.enable(TE_F3D5PHI3X1_F4D5PHI2X1_SP_F3D5PHI3X1_F4D5PHI2X1_wr_en),
.number_out(SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5),
.start(TE_F3D5PHI3X1_F4D5PHI2X1_start),
.done(SP_F3D5PHI3X1_F4D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI3X1_F4D5PHI3X1_SP_F3D5PHI3X1_F4D5PHI3X1;
wire TE_F3D5PHI3X1_F4D5PHI3X1_SP_F3D5PHI3X1_F4D5PHI3X1_wr_en;
wire [5:0] SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI3X1_F4D5PHI3X1(
.data_in(TE_F3D5PHI3X1_F4D5PHI3X1_SP_F3D5PHI3X1_F4D5PHI3X1),
.enable(TE_F3D5PHI3X1_F4D5PHI3X1_SP_F3D5PHI3X1_F4D5PHI3X1_wr_en),
.number_out(SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5),
.start(TE_F3D5PHI3X1_F4D5PHI3X1_start),
.done(SP_F3D5PHI3X1_F4D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI4X1_F4D5PHI3X1_SP_F3D5PHI4X1_F4D5PHI3X1;
wire TE_F3D5PHI4X1_F4D5PHI3X1_SP_F3D5PHI4X1_F4D5PHI3X1_wr_en;
wire [5:0] SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI4X1_F4D5PHI3X1(
.data_in(TE_F3D5PHI4X1_F4D5PHI3X1_SP_F3D5PHI4X1_F4D5PHI3X1),
.enable(TE_F3D5PHI4X1_F4D5PHI3X1_SP_F3D5PHI4X1_F4D5PHI3X1_wr_en),
.number_out(SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5),
.start(TE_F3D5PHI4X1_F4D5PHI3X1_start),
.done(SP_F3D5PHI4X1_F4D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI1X1_F4D5PHI1X2_SP_F3D5PHI1X1_F4D5PHI1X2;
wire TE_F3D5PHI1X1_F4D5PHI1X2_SP_F3D5PHI1X1_F4D5PHI1X2_wr_en;
wire [5:0] SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI1X1_F4D5PHI1X2(
.data_in(TE_F3D5PHI1X1_F4D5PHI1X2_SP_F3D5PHI1X1_F4D5PHI1X2),
.enable(TE_F3D5PHI1X1_F4D5PHI1X2_SP_F3D5PHI1X1_F4D5PHI1X2_wr_en),
.number_out(SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5),
.start(TE_F3D5PHI1X1_F4D5PHI1X2_start),
.done(SP_F3D5PHI1X1_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI2X1_F4D5PHI1X2_SP_F3D5PHI2X1_F4D5PHI1X2;
wire TE_F3D5PHI2X1_F4D5PHI1X2_SP_F3D5PHI2X1_F4D5PHI1X2_wr_en;
wire [5:0] SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI2X1_F4D5PHI1X2(
.data_in(TE_F3D5PHI2X1_F4D5PHI1X2_SP_F3D5PHI2X1_F4D5PHI1X2),
.enable(TE_F3D5PHI2X1_F4D5PHI1X2_SP_F3D5PHI2X1_F4D5PHI1X2_wr_en),
.number_out(SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5),
.start(TE_F3D5PHI2X1_F4D5PHI1X2_start),
.done(SP_F3D5PHI2X1_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI2X1_F4D5PHI2X2_SP_F3D5PHI2X1_F4D5PHI2X2;
wire TE_F3D5PHI2X1_F4D5PHI2X2_SP_F3D5PHI2X1_F4D5PHI2X2_wr_en;
wire [5:0] SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI2X1_F4D5PHI2X2(
.data_in(TE_F3D5PHI2X1_F4D5PHI2X2_SP_F3D5PHI2X1_F4D5PHI2X2),
.enable(TE_F3D5PHI2X1_F4D5PHI2X2_SP_F3D5PHI2X1_F4D5PHI2X2_wr_en),
.number_out(SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5),
.start(TE_F3D5PHI2X1_F4D5PHI2X2_start),
.done(SP_F3D5PHI2X1_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI3X1_F4D5PHI2X2_SP_F3D5PHI3X1_F4D5PHI2X2;
wire TE_F3D5PHI3X1_F4D5PHI2X2_SP_F3D5PHI3X1_F4D5PHI2X2_wr_en;
wire [5:0] SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI3X1_F4D5PHI2X2(
.data_in(TE_F3D5PHI3X1_F4D5PHI2X2_SP_F3D5PHI3X1_F4D5PHI2X2),
.enable(TE_F3D5PHI3X1_F4D5PHI2X2_SP_F3D5PHI3X1_F4D5PHI2X2_wr_en),
.number_out(SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5),
.start(TE_F3D5PHI3X1_F4D5PHI2X2_start),
.done(SP_F3D5PHI3X1_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI3X1_F4D5PHI3X2_SP_F3D5PHI3X1_F4D5PHI3X2;
wire TE_F3D5PHI3X1_F4D5PHI3X2_SP_F3D5PHI3X1_F4D5PHI3X2_wr_en;
wire [5:0] SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI3X1_F4D5PHI3X2(
.data_in(TE_F3D5PHI3X1_F4D5PHI3X2_SP_F3D5PHI3X1_F4D5PHI3X2),
.enable(TE_F3D5PHI3X1_F4D5PHI3X2_SP_F3D5PHI3X1_F4D5PHI3X2_wr_en),
.number_out(SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5),
.start(TE_F3D5PHI3X1_F4D5PHI3X2_start),
.done(SP_F3D5PHI3X1_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI4X1_F4D5PHI3X2_SP_F3D5PHI4X1_F4D5PHI3X2;
wire TE_F3D5PHI4X1_F4D5PHI3X2_SP_F3D5PHI4X1_F4D5PHI3X2_wr_en;
wire [5:0] SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI4X1_F4D5PHI3X2(
.data_in(TE_F3D5PHI4X1_F4D5PHI3X2_SP_F3D5PHI4X1_F4D5PHI3X2),
.enable(TE_F3D5PHI4X1_F4D5PHI3X2_SP_F3D5PHI4X1_F4D5PHI3X2_wr_en),
.number_out(SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5),
.start(TE_F3D5PHI4X1_F4D5PHI3X2_start),
.done(SP_F3D5PHI4X1_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI1X2_F4D5PHI1X2_SP_F3D5PHI1X2_F4D5PHI1X2;
wire TE_F3D5PHI1X2_F4D5PHI1X2_SP_F3D5PHI1X2_F4D5PHI1X2_wr_en;
wire [5:0] SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI1X2_F4D5PHI1X2(
.data_in(TE_F3D5PHI1X2_F4D5PHI1X2_SP_F3D5PHI1X2_F4D5PHI1X2),
.enable(TE_F3D5PHI1X2_F4D5PHI1X2_SP_F3D5PHI1X2_F4D5PHI1X2_wr_en),
.number_out(SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5),
.start(TE_F3D5PHI1X2_F4D5PHI1X2_start),
.done(SP_F3D5PHI1X2_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI2X2_F4D5PHI1X2_SP_F3D5PHI2X2_F4D5PHI1X2;
wire TE_F3D5PHI2X2_F4D5PHI1X2_SP_F3D5PHI2X2_F4D5PHI1X2_wr_en;
wire [5:0] SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI2X2_F4D5PHI1X2(
.data_in(TE_F3D5PHI2X2_F4D5PHI1X2_SP_F3D5PHI2X2_F4D5PHI1X2),
.enable(TE_F3D5PHI2X2_F4D5PHI1X2_SP_F3D5PHI2X2_F4D5PHI1X2_wr_en),
.number_out(SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5),
.start(TE_F3D5PHI2X2_F4D5PHI1X2_start),
.done(SP_F3D5PHI2X2_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI2X2_F4D5PHI2X2_SP_F3D5PHI2X2_F4D5PHI2X2;
wire TE_F3D5PHI2X2_F4D5PHI2X2_SP_F3D5PHI2X2_F4D5PHI2X2_wr_en;
wire [5:0] SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI2X2_F4D5PHI2X2(
.data_in(TE_F3D5PHI2X2_F4D5PHI2X2_SP_F3D5PHI2X2_F4D5PHI2X2),
.enable(TE_F3D5PHI2X2_F4D5PHI2X2_SP_F3D5PHI2X2_F4D5PHI2X2_wr_en),
.number_out(SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5),
.start(TE_F3D5PHI2X2_F4D5PHI2X2_start),
.done(SP_F3D5PHI2X2_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI3X2_F4D5PHI2X2_SP_F3D5PHI3X2_F4D5PHI2X2;
wire TE_F3D5PHI3X2_F4D5PHI2X2_SP_F3D5PHI3X2_F4D5PHI2X2_wr_en;
wire [5:0] SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI3X2_F4D5PHI2X2(
.data_in(TE_F3D5PHI3X2_F4D5PHI2X2_SP_F3D5PHI3X2_F4D5PHI2X2),
.enable(TE_F3D5PHI3X2_F4D5PHI2X2_SP_F3D5PHI3X2_F4D5PHI2X2_wr_en),
.number_out(SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5),
.start(TE_F3D5PHI3X2_F4D5PHI2X2_start),
.done(SP_F3D5PHI3X2_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI3X2_F4D5PHI3X2_SP_F3D5PHI3X2_F4D5PHI3X2;
wire TE_F3D5PHI3X2_F4D5PHI3X2_SP_F3D5PHI3X2_F4D5PHI3X2_wr_en;
wire [5:0] SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI3X2_F4D5PHI3X2(
.data_in(TE_F3D5PHI3X2_F4D5PHI3X2_SP_F3D5PHI3X2_F4D5PHI3X2),
.enable(TE_F3D5PHI3X2_F4D5PHI3X2_SP_F3D5PHI3X2_F4D5PHI3X2_wr_en),
.number_out(SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5),
.start(TE_F3D5PHI3X2_F4D5PHI3X2_start),
.done(SP_F3D5PHI3X2_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_F3D5PHI4X2_F4D5PHI3X2_SP_F3D5PHI4X2_F4D5PHI3X2;
wire TE_F3D5PHI4X2_F4D5PHI3X2_SP_F3D5PHI4X2_F4D5PHI3X2_wr_en;
wire [5:0] SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5_number;
wire [8:0] SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5_read_add;
wire [11:0] SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5;
StubPairs  SP_F3D5PHI4X2_F4D5PHI3X2(
.data_in(TE_F3D5PHI4X2_F4D5PHI3X2_SP_F3D5PHI4X2_F4D5PHI3X2),
.enable(TE_F3D5PHI4X2_F4D5PHI3X2_SP_F3D5PHI4X2_F4D5PHI3X2_wr_en),
.number_out(SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5_number),
.read_add(SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5_read_add),
.data_out(SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5),
.start(TE_F3D5PHI4X2_F4D5PHI3X2_start),
.done(SP_F3D5PHI4X2_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F3D5_AS_F3D5n1;
wire VMRD_F3D5_AS_F3D5n1_wr_en;
wire [10:0] AS_F3D5n1_TC_F3D5F4D5_read_add;
wire [35:0] AS_F3D5n1_TC_F3D5F4D5;
AllStubs  AS_F3D5n1(
.data_in(VMRD_F3D5_AS_F3D5n1),
.enable(VMRD_F3D5_AS_F3D5n1_wr_en),
.read_add(AS_F3D5n1_TC_F3D5F4D5_read_add),
.data_out(AS_F3D5n1_TC_F3D5F4D5),
.start(VMRD_F3D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F4D5_AS_F4D5n1;
wire VMRD_F4D5_AS_F4D5n1_wr_en;
wire [10:0] AS_F4D5n1_TC_F3D5F4D5_read_add;
wire [35:0] AS_F4D5n1_TC_F3D5F4D5;
AllStubs  AS_F4D5n1(
.data_in(VMRD_F4D5_AS_F4D5n1),
.enable(VMRD_F4D5_AS_F4D5n1_wr_en),
.read_add(AS_F4D5n1_TC_F3D5F4D5_read_add),
.data_out(AS_F4D5n1_TC_F3D5F4D5),
.start(VMRD_F4D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Plus_TPROJ_FromPlus_F3D5_F1F2;
wire PT_L3F3F5_Plus_TPROJ_FromPlus_F3D5_F1F2_wr_en;
wire [5:0] TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2_number;
wire [9:0] TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2_read_add;
wire [53:0] TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2;
TrackletProjections #(1'b1) TPROJ_FromPlus_F3D5_F1F2(
.data_in(PT_L3F3F5_Plus_TPROJ_FromPlus_F3D5_F1F2),
.enable(PT_L3F3F5_Plus_TPROJ_FromPlus_F3D5_F1F2_wr_en),
.number_out(TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2_number),
.read_add(TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2_read_add),
.data_out(TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2),
.start(PT_L3F3F5_Plus_start),
.done(TPROJ_FromPlus_F3D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Minus_TPROJ_FromMinus_F3D5_F1F2;
wire PT_L3F3F5_Minus_TPROJ_FromMinus_F3D5_F1F2_wr_en;
wire [5:0] TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2_number;
wire [9:0] TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2_read_add;
wire [53:0] TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2;
TrackletProjections #(1'b1) TPROJ_FromMinus_F3D5_F1F2(
.data_in(PT_L3F3F5_Minus_TPROJ_FromMinus_F3D5_F1F2),
.enable(PT_L3F3F5_Minus_TPROJ_FromMinus_F3D5_F1F2_wr_en),
.number_out(TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2_number),
.read_add(TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2_read_add),
.data_out(TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2),
.start(PT_L3F3F5_Minus_start),
.done(TPROJ_FromMinus_F3D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F1D5F2D5_TPROJ_F1D5F2D5_F3D5;
wire TC_F1D5F2D5_TPROJ_F1D5F2D5_F3D5_wr_en;
wire [5:0] TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2_number;
wire [9:0] TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2_read_add;
wire [53:0] TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2;
TrackletProjections  TPROJ_F1D5F2D5_F3D5(
.data_in(TC_F1D5F2D5_TPROJ_F1D5F2D5_F3D5),
.enable(TC_F1D5F2D5_TPROJ_F1D5F2D5_F3D5_wr_en),
.number_out(TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2_number),
.read_add(TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2_read_add),
.data_out(TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_F1D5F2D5_F3D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_F4D5_F1F2;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_F4D5_F1F2_wr_en;
wire [5:0] TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2_number;
wire [9:0] TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2_read_add;
wire [53:0] TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2;
TrackletProjections #(1'b1) TPROJ_FromPlus_F4D5_F1F2(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_F4D5_F1F2),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_F4D5_F1F2_wr_en),
.number_out(TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2_number),
.read_add(TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2_read_add),
.data_out(TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_F4D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_F4D5_F1F2;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_F4D5_F1F2_wr_en;
wire [5:0] TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2_number;
wire [9:0] TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2_read_add;
wire [53:0] TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2;
TrackletProjections #(1'b1) TPROJ_FromMinus_F4D5_F1F2(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_F4D5_F1F2),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_F4D5_F1F2_wr_en),
.number_out(TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2_number),
.read_add(TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2_read_add),
.data_out(TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_F4D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F1D5F2D5_TPROJ_F1D5F2D5_F4D5;
wire TC_F1D5F2D5_TPROJ_F1D5F2D5_F4D5_wr_en;
wire [5:0] TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2_number;
wire [9:0] TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2_read_add;
wire [53:0] TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2;
TrackletProjections  TPROJ_F1D5F2D5_F4D5(
.data_in(TC_F1D5F2D5_TPROJ_F1D5F2D5_F4D5),
.enable(TC_F1D5F2D5_TPROJ_F1D5F2D5_F4D5_wr_en),
.number_out(TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2_number),
.read_add(TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2_read_add),
.data_out(TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_F1D5F2D5_F4D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F1F2;
wire PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F1F2_wr_en;
wire [5:0] TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2_number;
wire [9:0] TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2_read_add;
wire [53:0] TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2;
TrackletProjections #(1'b1) TPROJ_FromPlus_F5D5_F1F2(
.data_in(PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F1F2),
.enable(PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F1F2_wr_en),
.number_out(TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2_number),
.read_add(TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2_read_add),
.data_out(TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2),
.start(PT_L3F3F5_Plus_start),
.done(TPROJ_FromPlus_F5D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F1F2;
wire PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F1F2_wr_en;
wire [5:0] TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2_number;
wire [9:0] TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2_read_add;
wire [53:0] TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2;
TrackletProjections #(1'b1) TPROJ_FromMinus_F5D5_F1F2(
.data_in(PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F1F2),
.enable(PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F1F2_wr_en),
.number_out(TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2_number),
.read_add(TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2_read_add),
.data_out(TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2),
.start(PT_L3F3F5_Minus_start),
.done(TPROJ_FromMinus_F5D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F1D5F2D5_TPROJ_F1D5F2D5_F5D5;
wire TC_F1D5F2D5_TPROJ_F1D5F2D5_F5D5_wr_en;
wire [5:0] TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2_number;
wire [9:0] TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2_read_add;
wire [53:0] TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2;
TrackletProjections  TPROJ_F1D5F2D5_F5D5(
.data_in(TC_F1D5F2D5_TPROJ_F1D5F2D5_F5D5),
.enable(TC_F1D5F2D5_TPROJ_F1D5F2D5_F5D5_wr_en),
.number_out(TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2_number),
.read_add(TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2_read_add),
.data_out(TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2),
.start(TC_F1D5F2D5_proj_start),
.done(TPROJ_F1D5F2D5_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Plus_TPROJ_FromPlus_F1D5_F3F4;
wire PT_F1L5_Plus_TPROJ_FromPlus_F1D5_F3F4_wr_en;
wire [5:0] TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4_number;
wire [9:0] TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4_read_add;
wire [53:0] TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4;
TrackletProjections #(1'b1) TPROJ_FromPlus_F1D5_F3F4(
.data_in(PT_F1L5_Plus_TPROJ_FromPlus_F1D5_F3F4),
.enable(PT_F1L5_Plus_TPROJ_FromPlus_F1D5_F3F4_wr_en),
.number_out(TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4_number),
.read_add(TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4_read_add),
.data_out(TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4),
.start(PT_F1L5_Plus_start),
.done(TPROJ_FromPlus_F1D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Minus_TPROJ_FromMinus_F1D5_F3F4;
wire PT_F1L5_Minus_TPROJ_FromMinus_F1D5_F3F4_wr_en;
wire [5:0] TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4_number;
wire [9:0] TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4_read_add;
wire [53:0] TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4;
TrackletProjections #(1'b1) TPROJ_FromMinus_F1D5_F3F4(
.data_in(PT_F1L5_Minus_TPROJ_FromMinus_F1D5_F3F4),
.enable(PT_F1L5_Minus_TPROJ_FromMinus_F1D5_F3F4_wr_en),
.number_out(TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4_number),
.read_add(TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4_read_add),
.data_out(TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4),
.start(PT_F1L5_Minus_start),
.done(TPROJ_FromMinus_F1D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_F3D5F4D5_F1D5;
wire TC_F3D5F4D5_TPROJ_F3D5F4D5_F1D5_wr_en;
wire [5:0] TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4_number;
wire [9:0] TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4_read_add;
wire [53:0] TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4;
TrackletProjections  TPROJ_F3D5F4D5_F1D5(
.data_in(TC_F3D5F4D5_TPROJ_F3D5F4D5_F1D5),
.enable(TC_F3D5F4D5_TPROJ_F3D5F4D5_F1D5_wr_en),
.number_out(TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4_number),
.read_add(TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4_read_add),
.data_out(TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_F3D5F4D5_F1D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_F2D5_F3F4;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_F2D5_F3F4_wr_en;
wire [5:0] TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4_number;
wire [9:0] TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4_read_add;
wire [53:0] TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4;
TrackletProjections #(1'b1) TPROJ_FromPlus_F2D5_F3F4(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_F2D5_F3F4),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_F2D5_F3F4_wr_en),
.number_out(TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4_number),
.read_add(TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4_read_add),
.data_out(TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_F2D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_F2D5_F3F4;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_F2D5_F3F4_wr_en;
wire [5:0] TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4_number;
wire [9:0] TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4_read_add;
wire [53:0] TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4;
TrackletProjections #(1'b1) TPROJ_FromMinus_F2D5_F3F4(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_F2D5_F3F4),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_F2D5_F3F4_wr_en),
.number_out(TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4_number),
.read_add(TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4_read_add),
.data_out(TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_F2D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_F3D5F4D5_F2D5;
wire TC_F3D5F4D5_TPROJ_F3D5F4D5_F2D5_wr_en;
wire [5:0] TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4_number;
wire [9:0] TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4_read_add;
wire [53:0] TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4;
TrackletProjections  TPROJ_F3D5F4D5_F2D5(
.data_in(TC_F3D5F4D5_TPROJ_F3D5F4D5_F2D5),
.enable(TC_F3D5F4D5_TPROJ_F3D5F4D5_F2D5_wr_en),
.number_out(TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4_number),
.read_add(TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4_read_add),
.data_out(TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_F3D5F4D5_F2D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F3F4;
wire PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F3F4_wr_en;
wire [5:0] TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4_number;
wire [9:0] TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4_read_add;
wire [53:0] TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4;
TrackletProjections #(1'b1) TPROJ_FromPlus_F5D5_F3F4(
.data_in(PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F3F4),
.enable(PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F3F4_wr_en),
.number_out(TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4_number),
.read_add(TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4_read_add),
.data_out(TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4),
.start(PT_L3F3F5_Plus_start),
.done(TPROJ_FromPlus_F5D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F3F4;
wire PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F3F4_wr_en;
wire [5:0] TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4_number;
wire [9:0] TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4_read_add;
wire [53:0] TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4;
TrackletProjections #(1'b1) TPROJ_FromMinus_F5D5_F3F4(
.data_in(PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F3F4),
.enable(PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F3F4_wr_en),
.number_out(TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4_number),
.read_add(TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4_read_add),
.data_out(TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4),
.start(PT_L3F3F5_Minus_start),
.done(TPROJ_FromMinus_F5D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_F3D5F4D5_TPROJ_F3D5F4D5_F5D5;
wire TC_F3D5F4D5_TPROJ_F3D5F4D5_F5D5_wr_en;
wire [5:0] TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4_number;
wire [9:0] TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4_read_add;
wire [53:0] TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4;
TrackletProjections  TPROJ_F3D5F4D5_F5D5(
.data_in(TC_F3D5F4D5_TPROJ_F3D5F4D5_F5D5),
.enable(TC_F3D5F4D5_TPROJ_F3D5F4D5_F5D5_wr_en),
.number_out(TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4_number),
.read_add(TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4_read_add),
.data_out(TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4),
.start(TC_F3D5F4D5_proj_start),
.done(TPROJ_F3D5F4D5_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X1;
wire PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X1_wr_en;
wire [5:0] VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1_number;
wire [8:0] VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1_read_add;
wire [13:0] VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1;
VMProjections  VMPROJ_F1F2_F3D5PHI1X1(
.data_in(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X1),
.enable(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X1_wr_en),
.number_out(VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1_number),
.read_add(VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1_read_add),
.data_out(VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1),
.start(PRD_F3D5_F1F2_start),
.done(VMPROJ_F1F2_F3D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI1X1n3;
wire VMRD_F3D5_VMS_F3D5PHI1X1n3_wr_en;
wire [5:0] VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1_number;
wire [10:0] VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1_read_add;
wire [18:0] VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1;
VMStubs #("Match") VMS_F3D5PHI1X1n3(
.data_in(VMRD_F3D5_VMS_F3D5PHI1X1n3),
.enable(VMRD_F3D5_VMS_F3D5PHI1X1n3_wr_en),
.number_out(VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1_number),
.read_add(VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1_read_add),
.data_out(VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X2;
wire PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X2_wr_en;
wire [5:0] VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2_number;
wire [8:0] VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2_read_add;
wire [13:0] VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2;
VMProjections  VMPROJ_F1F2_F3D5PHI1X2(
.data_in(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X2),
.enable(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X2_wr_en),
.number_out(VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2_number),
.read_add(VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2_read_add),
.data_out(VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2),
.start(PRD_F3D5_F1F2_start),
.done(VMPROJ_F1F2_F3D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI1X2n2;
wire VMRD_F3D5_VMS_F3D5PHI1X2n2_wr_en;
wire [5:0] VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2_number;
wire [10:0] VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2_read_add;
wire [18:0] VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2;
VMStubs #("Match") VMS_F3D5PHI1X2n2(
.data_in(VMRD_F3D5_VMS_F3D5PHI1X2n2),
.enable(VMRD_F3D5_VMS_F3D5PHI1X2n2_wr_en),
.number_out(VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2_number),
.read_add(VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2_read_add),
.data_out(VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X1;
wire PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X1_wr_en;
wire [5:0] VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1_number;
wire [8:0] VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1_read_add;
wire [13:0] VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1;
VMProjections  VMPROJ_F1F2_F3D5PHI2X1(
.data_in(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X1),
.enable(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X1_wr_en),
.number_out(VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1_number),
.read_add(VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1_read_add),
.data_out(VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1),
.start(PRD_F3D5_F1F2_start),
.done(VMPROJ_F1F2_F3D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI2X1n5;
wire VMRD_F3D5_VMS_F3D5PHI2X1n5_wr_en;
wire [5:0] VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1_number;
wire [10:0] VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1_read_add;
wire [18:0] VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1;
VMStubs #("Match") VMS_F3D5PHI2X1n5(
.data_in(VMRD_F3D5_VMS_F3D5PHI2X1n5),
.enable(VMRD_F3D5_VMS_F3D5PHI2X1n5_wr_en),
.number_out(VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1_number),
.read_add(VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1_read_add),
.data_out(VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X2;
wire PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X2_wr_en;
wire [5:0] VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2_number;
wire [8:0] VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2_read_add;
wire [13:0] VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2;
VMProjections  VMPROJ_F1F2_F3D5PHI2X2(
.data_in(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X2),
.enable(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X2_wr_en),
.number_out(VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2_number),
.read_add(VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2_read_add),
.data_out(VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2),
.start(PRD_F3D5_F1F2_start),
.done(VMPROJ_F1F2_F3D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI2X2n3;
wire VMRD_F3D5_VMS_F3D5PHI2X2n3_wr_en;
wire [5:0] VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2_number;
wire [10:0] VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2_read_add;
wire [18:0] VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2;
VMStubs #("Match") VMS_F3D5PHI2X2n3(
.data_in(VMRD_F3D5_VMS_F3D5PHI2X2n3),
.enable(VMRD_F3D5_VMS_F3D5PHI2X2n3_wr_en),
.number_out(VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2_number),
.read_add(VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2_read_add),
.data_out(VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X1;
wire PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X1_wr_en;
wire [5:0] VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1_number;
wire [8:0] VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1_read_add;
wire [13:0] VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1;
VMProjections  VMPROJ_F1F2_F3D5PHI3X1(
.data_in(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X1),
.enable(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X1_wr_en),
.number_out(VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1_number),
.read_add(VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1_read_add),
.data_out(VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1),
.start(PRD_F3D5_F1F2_start),
.done(VMPROJ_F1F2_F3D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI3X1n5;
wire VMRD_F3D5_VMS_F3D5PHI3X1n5_wr_en;
wire [5:0] VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1_number;
wire [10:0] VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1_read_add;
wire [18:0] VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1;
VMStubs #("Match") VMS_F3D5PHI3X1n5(
.data_in(VMRD_F3D5_VMS_F3D5PHI3X1n5),
.enable(VMRD_F3D5_VMS_F3D5PHI3X1n5_wr_en),
.number_out(VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1_number),
.read_add(VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1_read_add),
.data_out(VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X2;
wire PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X2_wr_en;
wire [5:0] VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2_number;
wire [8:0] VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2_read_add;
wire [13:0] VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2;
VMProjections  VMPROJ_F1F2_F3D5PHI3X2(
.data_in(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X2),
.enable(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X2_wr_en),
.number_out(VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2_number),
.read_add(VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2_read_add),
.data_out(VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2),
.start(PRD_F3D5_F1F2_start),
.done(VMPROJ_F1F2_F3D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI3X2n3;
wire VMRD_F3D5_VMS_F3D5PHI3X2n3_wr_en;
wire [5:0] VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2_number;
wire [10:0] VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2_read_add;
wire [18:0] VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2;
VMStubs #("Match") VMS_F3D5PHI3X2n3(
.data_in(VMRD_F3D5_VMS_F3D5PHI3X2n3),
.enable(VMRD_F3D5_VMS_F3D5PHI3X2n3_wr_en),
.number_out(VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2_number),
.read_add(VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2_read_add),
.data_out(VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X1;
wire PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X1_wr_en;
wire [5:0] VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1_number;
wire [8:0] VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1_read_add;
wire [13:0] VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1;
VMProjections  VMPROJ_F1F2_F3D5PHI4X1(
.data_in(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X1),
.enable(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X1_wr_en),
.number_out(VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1_number),
.read_add(VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1_read_add),
.data_out(VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1),
.start(PRD_F3D5_F1F2_start),
.done(VMPROJ_F1F2_F3D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI4X1n3;
wire VMRD_F3D5_VMS_F3D5PHI4X1n3_wr_en;
wire [5:0] VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1_number;
wire [10:0] VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1_read_add;
wire [18:0] VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1;
VMStubs #("Match") VMS_F3D5PHI4X1n3(
.data_in(VMRD_F3D5_VMS_F3D5PHI4X1n3),
.enable(VMRD_F3D5_VMS_F3D5PHI4X1n3_wr_en),
.number_out(VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1_number),
.read_add(VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1_read_add),
.data_out(VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI4X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X2;
wire PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X2_wr_en;
wire [5:0] VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2_number;
wire [8:0] VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2_read_add;
wire [13:0] VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2;
VMProjections  VMPROJ_F1F2_F3D5PHI4X2(
.data_in(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X2),
.enable(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X2_wr_en),
.number_out(VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2_number),
.read_add(VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2_read_add),
.data_out(VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2),
.start(PRD_F3D5_F1F2_start),
.done(VMPROJ_F1F2_F3D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F3D5_VMS_F3D5PHI4X2n2;
wire VMRD_F3D5_VMS_F3D5PHI4X2n2_wr_en;
wire [5:0] VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2_number;
wire [10:0] VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2_read_add;
wire [18:0] VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2;
VMStubs #("Match") VMS_F3D5PHI4X2n2(
.data_in(VMRD_F3D5_VMS_F3D5PHI4X2n2),
.enable(VMRD_F3D5_VMS_F3D5PHI4X2n2_wr_en),
.number_out(VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2_number),
.read_add(VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2_read_add),
.data_out(VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2),
.start(VMRD_F3D5_start),
.done(VMS_F3D5PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X1;
wire PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X1_wr_en;
wire [5:0] VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1_number;
wire [8:0] VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1_read_add;
wire [13:0] VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1;
VMProjections  VMPROJ_F1F2_F4D5PHI1X1(
.data_in(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X1),
.enable(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X1_wr_en),
.number_out(VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1_number),
.read_add(VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1_read_add),
.data_out(VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1),
.start(PRD_F4D5_F1F2_start),
.done(VMPROJ_F1F2_F4D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI1X1n3;
wire VMRD_F4D5_VMS_F4D5PHI1X1n3_wr_en;
wire [5:0] VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1_number;
wire [10:0] VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1_read_add;
wire [18:0] VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1;
VMStubs #("Match") VMS_F4D5PHI1X1n3(
.data_in(VMRD_F4D5_VMS_F4D5PHI1X1n3),
.enable(VMRD_F4D5_VMS_F4D5PHI1X1n3_wr_en),
.number_out(VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1_number),
.read_add(VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1_read_add),
.data_out(VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X2;
wire PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X2_wr_en;
wire [5:0] VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2_number;
wire [8:0] VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2_read_add;
wire [13:0] VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2;
VMProjections  VMPROJ_F1F2_F4D5PHI1X2(
.data_in(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X2),
.enable(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X2_wr_en),
.number_out(VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2_number),
.read_add(VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2_read_add),
.data_out(VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2),
.start(PRD_F4D5_F1F2_start),
.done(VMPROJ_F1F2_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI1X2n5;
wire VMRD_F4D5_VMS_F4D5PHI1X2n5_wr_en;
wire [5:0] VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2_number;
wire [10:0] VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2_read_add;
wire [18:0] VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2;
VMStubs #("Match") VMS_F4D5PHI1X2n5(
.data_in(VMRD_F4D5_VMS_F4D5PHI1X2n5),
.enable(VMRD_F4D5_VMS_F4D5PHI1X2n5_wr_en),
.number_out(VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2_number),
.read_add(VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2_read_add),
.data_out(VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI1X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X1;
wire PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X1_wr_en;
wire [5:0] VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1_number;
wire [8:0] VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1_read_add;
wire [13:0] VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1;
VMProjections  VMPROJ_F1F2_F4D5PHI2X1(
.data_in(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X1),
.enable(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X1_wr_en),
.number_out(VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1_number),
.read_add(VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1_read_add),
.data_out(VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1),
.start(PRD_F4D5_F1F2_start),
.done(VMPROJ_F1F2_F4D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI2X1n3;
wire VMRD_F4D5_VMS_F4D5PHI2X1n3_wr_en;
wire [5:0] VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1_number;
wire [10:0] VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1_read_add;
wire [18:0] VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1;
VMStubs #("Match") VMS_F4D5PHI2X1n3(
.data_in(VMRD_F4D5_VMS_F4D5PHI2X1n3),
.enable(VMRD_F4D5_VMS_F4D5PHI2X1n3_wr_en),
.number_out(VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1_number),
.read_add(VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1_read_add),
.data_out(VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X2;
wire PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X2_wr_en;
wire [5:0] VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2_number;
wire [8:0] VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2_read_add;
wire [13:0] VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2;
VMProjections  VMPROJ_F1F2_F4D5PHI2X2(
.data_in(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X2),
.enable(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X2_wr_en),
.number_out(VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2_number),
.read_add(VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2_read_add),
.data_out(VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2),
.start(PRD_F4D5_F1F2_start),
.done(VMPROJ_F1F2_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI2X2n5;
wire VMRD_F4D5_VMS_F4D5PHI2X2n5_wr_en;
wire [5:0] VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2_number;
wire [10:0] VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2_read_add;
wire [18:0] VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2;
VMStubs #("Match") VMS_F4D5PHI2X2n5(
.data_in(VMRD_F4D5_VMS_F4D5PHI2X2n5),
.enable(VMRD_F4D5_VMS_F4D5PHI2X2n5_wr_en),
.number_out(VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2_number),
.read_add(VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2_read_add),
.data_out(VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X1;
wire PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X1_wr_en;
wire [5:0] VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1_number;
wire [8:0] VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1_read_add;
wire [13:0] VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1;
VMProjections  VMPROJ_F1F2_F4D5PHI3X1(
.data_in(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X1),
.enable(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X1_wr_en),
.number_out(VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1_number),
.read_add(VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1_read_add),
.data_out(VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1),
.start(PRD_F4D5_F1F2_start),
.done(VMPROJ_F1F2_F4D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI3X1n3;
wire VMRD_F4D5_VMS_F4D5PHI3X1n3_wr_en;
wire [5:0] VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1_number;
wire [10:0] VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1_read_add;
wire [18:0] VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1;
VMStubs #("Match") VMS_F4D5PHI3X1n3(
.data_in(VMRD_F4D5_VMS_F4D5PHI3X1n3),
.enable(VMRD_F4D5_VMS_F4D5PHI3X1n3_wr_en),
.number_out(VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1_number),
.read_add(VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1_read_add),
.data_out(VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X2;
wire PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X2_wr_en;
wire [5:0] VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2_number;
wire [8:0] VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2_read_add;
wire [13:0] VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2;
VMProjections  VMPROJ_F1F2_F4D5PHI3X2(
.data_in(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X2),
.enable(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X2_wr_en),
.number_out(VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2_number),
.read_add(VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2_read_add),
.data_out(VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2),
.start(PRD_F4D5_F1F2_start),
.done(VMPROJ_F1F2_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F4D5_VMS_F4D5PHI3X2n5;
wire VMRD_F4D5_VMS_F4D5PHI3X2n5_wr_en;
wire [5:0] VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2_number;
wire [10:0] VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2_read_add;
wire [18:0] VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2;
VMStubs #("Match") VMS_F4D5PHI3X2n5(
.data_in(VMRD_F4D5_VMS_F4D5PHI3X2n5),
.enable(VMRD_F4D5_VMS_F4D5PHI3X2n5_wr_en),
.number_out(VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2_number),
.read_add(VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2_read_add),
.data_out(VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2),
.start(VMRD_F4D5_start),
.done(VMS_F4D5PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X1;
wire PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X1_wr_en;
wire [5:0] VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1_number;
wire [8:0] VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1_read_add;
wire [13:0] VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1;
VMProjections  VMPROJ_F1F2_F5D5PHI1X1(
.data_in(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X1),
.enable(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X1_wr_en),
.number_out(VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1_number),
.read_add(VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1_read_add),
.data_out(VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1),
.start(PRD_F5D5_F1F2_start),
.done(VMPROJ_F1F2_F5D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI1X1n1;
wire VMRD_F5D5_VMS_F5D5PHI1X1n1_wr_en;
wire [5:0] VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1_number;
wire [10:0] VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1_read_add;
wire [18:0] VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1;
VMStubs #("Match") VMS_F5D5PHI1X1n1(
.data_in(VMRD_F5D5_VMS_F5D5PHI1X1n1),
.enable(VMRD_F5D5_VMS_F5D5PHI1X1n1_wr_en),
.number_out(VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1_number),
.read_add(VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1_read_add),
.data_out(VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X2;
wire PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X2_wr_en;
wire [5:0] VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2_number;
wire [8:0] VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2_read_add;
wire [13:0] VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2;
VMProjections  VMPROJ_F1F2_F5D5PHI1X2(
.data_in(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X2),
.enable(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X2_wr_en),
.number_out(VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2_number),
.read_add(VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2_read_add),
.data_out(VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2),
.start(PRD_F5D5_F1F2_start),
.done(VMPROJ_F1F2_F5D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI1X2n1;
wire VMRD_F5D5_VMS_F5D5PHI1X2n1_wr_en;
wire [5:0] VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2_number;
wire [10:0] VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2_read_add;
wire [18:0] VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2;
VMStubs #("Match") VMS_F5D5PHI1X2n1(
.data_in(VMRD_F5D5_VMS_F5D5PHI1X2n1),
.enable(VMRD_F5D5_VMS_F5D5PHI1X2n1_wr_en),
.number_out(VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2_number),
.read_add(VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2_read_add),
.data_out(VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X1;
wire PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X1_wr_en;
wire [5:0] VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1_number;
wire [8:0] VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1_read_add;
wire [13:0] VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1;
VMProjections  VMPROJ_F1F2_F5D5PHI2X1(
.data_in(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X1),
.enable(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X1_wr_en),
.number_out(VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1_number),
.read_add(VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1_read_add),
.data_out(VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1),
.start(PRD_F5D5_F1F2_start),
.done(VMPROJ_F1F2_F5D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI2X1n1;
wire VMRD_F5D5_VMS_F5D5PHI2X1n1_wr_en;
wire [5:0] VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1_number;
wire [10:0] VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1_read_add;
wire [18:0] VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1;
VMStubs #("Match") VMS_F5D5PHI2X1n1(
.data_in(VMRD_F5D5_VMS_F5D5PHI2X1n1),
.enable(VMRD_F5D5_VMS_F5D5PHI2X1n1_wr_en),
.number_out(VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1_number),
.read_add(VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1_read_add),
.data_out(VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X2;
wire PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X2_wr_en;
wire [5:0] VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2_number;
wire [8:0] VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2_read_add;
wire [13:0] VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2;
VMProjections  VMPROJ_F1F2_F5D5PHI2X2(
.data_in(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X2),
.enable(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X2_wr_en),
.number_out(VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2_number),
.read_add(VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2_read_add),
.data_out(VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2),
.start(PRD_F5D5_F1F2_start),
.done(VMPROJ_F1F2_F5D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI2X2n1;
wire VMRD_F5D5_VMS_F5D5PHI2X2n1_wr_en;
wire [5:0] VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2_number;
wire [10:0] VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2_read_add;
wire [18:0] VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2;
VMStubs #("Match") VMS_F5D5PHI2X2n1(
.data_in(VMRD_F5D5_VMS_F5D5PHI2X2n1),
.enable(VMRD_F5D5_VMS_F5D5PHI2X2n1_wr_en),
.number_out(VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2_number),
.read_add(VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2_read_add),
.data_out(VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X1;
wire PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X1_wr_en;
wire [5:0] VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1_number;
wire [8:0] VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1_read_add;
wire [13:0] VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1;
VMProjections  VMPROJ_F1F2_F5D5PHI3X1(
.data_in(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X1),
.enable(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X1_wr_en),
.number_out(VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1_number),
.read_add(VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1_read_add),
.data_out(VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1),
.start(PRD_F5D5_F1F2_start),
.done(VMPROJ_F1F2_F5D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI3X1n1;
wire VMRD_F5D5_VMS_F5D5PHI3X1n1_wr_en;
wire [5:0] VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1_number;
wire [10:0] VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1_read_add;
wire [18:0] VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1;
VMStubs #("Match") VMS_F5D5PHI3X1n1(
.data_in(VMRD_F5D5_VMS_F5D5PHI3X1n1),
.enable(VMRD_F5D5_VMS_F5D5PHI3X1n1_wr_en),
.number_out(VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1_number),
.read_add(VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1_read_add),
.data_out(VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X2;
wire PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X2_wr_en;
wire [5:0] VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2_number;
wire [8:0] VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2_read_add;
wire [13:0] VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2;
VMProjections  VMPROJ_F1F2_F5D5PHI3X2(
.data_in(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X2),
.enable(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X2_wr_en),
.number_out(VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2_number),
.read_add(VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2_read_add),
.data_out(VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2),
.start(PRD_F5D5_F1F2_start),
.done(VMPROJ_F1F2_F5D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI3X2n1;
wire VMRD_F5D5_VMS_F5D5PHI3X2n1_wr_en;
wire [5:0] VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2_number;
wire [10:0] VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2_read_add;
wire [18:0] VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2;
VMStubs #("Match") VMS_F5D5PHI3X2n1(
.data_in(VMRD_F5D5_VMS_F5D5PHI3X2n1),
.enable(VMRD_F5D5_VMS_F5D5PHI3X2n1_wr_en),
.number_out(VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2_number),
.read_add(VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2_read_add),
.data_out(VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X1;
wire PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X1_wr_en;
wire [5:0] VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1_number;
wire [8:0] VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1_read_add;
wire [13:0] VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1;
VMProjections  VMPROJ_F1F2_F5D5PHI4X1(
.data_in(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X1),
.enable(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X1_wr_en),
.number_out(VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1_number),
.read_add(VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1_read_add),
.data_out(VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1),
.start(PRD_F5D5_F1F2_start),
.done(VMPROJ_F1F2_F5D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI4X1n1;
wire VMRD_F5D5_VMS_F5D5PHI4X1n1_wr_en;
wire [5:0] VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1_number;
wire [10:0] VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1_read_add;
wire [18:0] VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1;
VMStubs #("Match") VMS_F5D5PHI4X1n1(
.data_in(VMRD_F5D5_VMS_F5D5PHI4X1n1),
.enable(VMRD_F5D5_VMS_F5D5PHI4X1n1_wr_en),
.number_out(VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1_number),
.read_add(VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1_read_add),
.data_out(VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X2;
wire PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X2_wr_en;
wire [5:0] VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2_number;
wire [8:0] VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2_read_add;
wire [13:0] VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2;
VMProjections  VMPROJ_F1F2_F5D5PHI4X2(
.data_in(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X2),
.enable(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X2_wr_en),
.number_out(VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2_number),
.read_add(VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2_read_add),
.data_out(VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2),
.start(PRD_F5D5_F1F2_start),
.done(VMPROJ_F1F2_F5D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI4X2n1;
wire VMRD_F5D5_VMS_F5D5PHI4X2n1_wr_en;
wire [5:0] VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2_number;
wire [10:0] VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2_read_add;
wire [18:0] VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2;
VMStubs #("Match") VMS_F5D5PHI4X2n1(
.data_in(VMRD_F5D5_VMS_F5D5PHI4X2n1),
.enable(VMRD_F5D5_VMS_F5D5PHI4X2n1_wr_en),
.number_out(VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2_number),
.read_add(VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2_read_add),
.data_out(VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X1;
wire PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X1_wr_en;
wire [5:0] VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1_number;
wire [8:0] VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1_read_add;
wire [13:0] VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1;
VMProjections  VMPROJ_F3F4_F1D5PHI1X1(
.data_in(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X1),
.enable(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X1_wr_en),
.number_out(VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1_number),
.read_add(VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1_read_add),
.data_out(VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1),
.start(PRD_F1D5_F3F4_start),
.done(VMPROJ_F3F4_F1D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI1X1n3;
wire VMRD_F1D5_VMS_F1D5PHI1X1n3_wr_en;
wire [5:0] VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1_number;
wire [10:0] VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1_read_add;
wire [18:0] VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1;
VMStubs #("Match") VMS_F1D5PHI1X1n3(
.data_in(VMRD_F1D5_VMS_F1D5PHI1X1n3),
.enable(VMRD_F1D5_VMS_F1D5PHI1X1n3_wr_en),
.number_out(VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1_number),
.read_add(VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1_read_add),
.data_out(VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X2;
wire PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X2_wr_en;
wire [5:0] VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2_number;
wire [8:0] VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2_read_add;
wire [13:0] VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2;
VMProjections  VMPROJ_F3F4_F1D5PHI1X2(
.data_in(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X2),
.enable(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X2_wr_en),
.number_out(VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2_number),
.read_add(VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2_read_add),
.data_out(VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2),
.start(PRD_F1D5_F3F4_start),
.done(VMPROJ_F3F4_F1D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI1X2n2;
wire VMRD_F1D5_VMS_F1D5PHI1X2n2_wr_en;
wire [5:0] VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2_number;
wire [10:0] VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2_read_add;
wire [18:0] VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2;
VMStubs #("Match") VMS_F1D5PHI1X2n2(
.data_in(VMRD_F1D5_VMS_F1D5PHI1X2n2),
.enable(VMRD_F1D5_VMS_F1D5PHI1X2n2_wr_en),
.number_out(VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2_number),
.read_add(VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2_read_add),
.data_out(VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X1;
wire PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X1_wr_en;
wire [5:0] VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1_number;
wire [8:0] VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1_read_add;
wire [13:0] VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1;
VMProjections  VMPROJ_F3F4_F1D5PHI2X1(
.data_in(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X1),
.enable(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X1_wr_en),
.number_out(VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1_number),
.read_add(VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1_read_add),
.data_out(VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1),
.start(PRD_F1D5_F3F4_start),
.done(VMPROJ_F3F4_F1D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI2X1n5;
wire VMRD_F1D5_VMS_F1D5PHI2X1n5_wr_en;
wire [5:0] VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1_number;
wire [10:0] VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1_read_add;
wire [18:0] VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1;
VMStubs #("Match") VMS_F1D5PHI2X1n5(
.data_in(VMRD_F1D5_VMS_F1D5PHI2X1n5),
.enable(VMRD_F1D5_VMS_F1D5PHI2X1n5_wr_en),
.number_out(VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1_number),
.read_add(VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1_read_add),
.data_out(VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X2;
wire PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X2_wr_en;
wire [5:0] VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2_number;
wire [8:0] VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2_read_add;
wire [13:0] VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2;
VMProjections  VMPROJ_F3F4_F1D5PHI2X2(
.data_in(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X2),
.enable(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X2_wr_en),
.number_out(VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2_number),
.read_add(VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2_read_add),
.data_out(VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2),
.start(PRD_F1D5_F3F4_start),
.done(VMPROJ_F3F4_F1D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI2X2n3;
wire VMRD_F1D5_VMS_F1D5PHI2X2n3_wr_en;
wire [5:0] VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2_number;
wire [10:0] VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2_read_add;
wire [18:0] VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2;
VMStubs #("Match") VMS_F1D5PHI2X2n3(
.data_in(VMRD_F1D5_VMS_F1D5PHI2X2n3),
.enable(VMRD_F1D5_VMS_F1D5PHI2X2n3_wr_en),
.number_out(VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2_number),
.read_add(VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2_read_add),
.data_out(VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X1;
wire PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X1_wr_en;
wire [5:0] VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1_number;
wire [8:0] VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1_read_add;
wire [13:0] VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1;
VMProjections  VMPROJ_F3F4_F1D5PHI3X1(
.data_in(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X1),
.enable(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X1_wr_en),
.number_out(VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1_number),
.read_add(VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1_read_add),
.data_out(VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1),
.start(PRD_F1D5_F3F4_start),
.done(VMPROJ_F3F4_F1D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI3X1n5;
wire VMRD_F1D5_VMS_F1D5PHI3X1n5_wr_en;
wire [5:0] VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1_number;
wire [10:0] VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1_read_add;
wire [18:0] VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1;
VMStubs #("Match") VMS_F1D5PHI3X1n5(
.data_in(VMRD_F1D5_VMS_F1D5PHI3X1n5),
.enable(VMRD_F1D5_VMS_F1D5PHI3X1n5_wr_en),
.number_out(VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1_number),
.read_add(VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1_read_add),
.data_out(VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X2;
wire PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X2_wr_en;
wire [5:0] VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2_number;
wire [8:0] VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2_read_add;
wire [13:0] VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2;
VMProjections  VMPROJ_F3F4_F1D5PHI3X2(
.data_in(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X2),
.enable(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X2_wr_en),
.number_out(VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2_number),
.read_add(VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2_read_add),
.data_out(VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2),
.start(PRD_F1D5_F3F4_start),
.done(VMPROJ_F3F4_F1D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI3X2n3;
wire VMRD_F1D5_VMS_F1D5PHI3X2n3_wr_en;
wire [5:0] VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2_number;
wire [10:0] VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2_read_add;
wire [18:0] VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2;
VMStubs #("Match") VMS_F1D5PHI3X2n3(
.data_in(VMRD_F1D5_VMS_F1D5PHI3X2n3),
.enable(VMRD_F1D5_VMS_F1D5PHI3X2n3_wr_en),
.number_out(VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2_number),
.read_add(VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2_read_add),
.data_out(VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X1;
wire PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X1_wr_en;
wire [5:0] VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1_number;
wire [8:0] VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1_read_add;
wire [13:0] VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1;
VMProjections  VMPROJ_F3F4_F1D5PHI4X1(
.data_in(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X1),
.enable(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X1_wr_en),
.number_out(VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1_number),
.read_add(VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1_read_add),
.data_out(VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1),
.start(PRD_F1D5_F3F4_start),
.done(VMPROJ_F3F4_F1D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI4X1n3;
wire VMRD_F1D5_VMS_F1D5PHI4X1n3_wr_en;
wire [5:0] VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1_number;
wire [10:0] VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1_read_add;
wire [18:0] VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1;
VMStubs #("Match") VMS_F1D5PHI4X1n3(
.data_in(VMRD_F1D5_VMS_F1D5PHI4X1n3),
.enable(VMRD_F1D5_VMS_F1D5PHI4X1n3_wr_en),
.number_out(VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1_number),
.read_add(VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1_read_add),
.data_out(VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI4X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X2;
wire PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X2_wr_en;
wire [5:0] VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2_number;
wire [8:0] VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2_read_add;
wire [13:0] VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2;
VMProjections  VMPROJ_F3F4_F1D5PHI4X2(
.data_in(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X2),
.enable(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X2_wr_en),
.number_out(VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2_number),
.read_add(VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2_read_add),
.data_out(VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2),
.start(PRD_F1D5_F3F4_start),
.done(VMPROJ_F3F4_F1D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F1D5_VMS_F1D5PHI4X2n2;
wire VMRD_F1D5_VMS_F1D5PHI4X2n2_wr_en;
wire [5:0] VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2_number;
wire [10:0] VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2_read_add;
wire [18:0] VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2;
VMStubs #("Match") VMS_F1D5PHI4X2n2(
.data_in(VMRD_F1D5_VMS_F1D5PHI4X2n2),
.enable(VMRD_F1D5_VMS_F1D5PHI4X2n2_wr_en),
.number_out(VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2_number),
.read_add(VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2_read_add),
.data_out(VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2),
.start(VMRD_F1D5_start),
.done(VMS_F1D5PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X1;
wire PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X1_wr_en;
wire [5:0] VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1_number;
wire [8:0] VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1_read_add;
wire [13:0] VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1;
VMProjections  VMPROJ_F3F4_F2D5PHI1X1(
.data_in(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X1),
.enable(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X1_wr_en),
.number_out(VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1_number),
.read_add(VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1_read_add),
.data_out(VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1),
.start(PRD_F2D5_F3F4_start),
.done(VMPROJ_F3F4_F2D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI1X1n3;
wire VMRD_F2D5_VMS_F2D5PHI1X1n3_wr_en;
wire [5:0] VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1_number;
wire [10:0] VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1_read_add;
wire [18:0] VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1;
VMStubs #("Match") VMS_F2D5PHI1X1n3(
.data_in(VMRD_F2D5_VMS_F2D5PHI1X1n3),
.enable(VMRD_F2D5_VMS_F2D5PHI1X1n3_wr_en),
.number_out(VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1_number),
.read_add(VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1_read_add),
.data_out(VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X2;
wire PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X2_wr_en;
wire [5:0] VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2_number;
wire [8:0] VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2_read_add;
wire [13:0] VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2;
VMProjections  VMPROJ_F3F4_F2D5PHI1X2(
.data_in(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X2),
.enable(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X2_wr_en),
.number_out(VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2_number),
.read_add(VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2_read_add),
.data_out(VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2),
.start(PRD_F2D5_F3F4_start),
.done(VMPROJ_F3F4_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI1X2n5;
wire VMRD_F2D5_VMS_F2D5PHI1X2n5_wr_en;
wire [5:0] VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2_number;
wire [10:0] VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2_read_add;
wire [18:0] VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2;
VMStubs #("Match") VMS_F2D5PHI1X2n5(
.data_in(VMRD_F2D5_VMS_F2D5PHI1X2n5),
.enable(VMRD_F2D5_VMS_F2D5PHI1X2n5_wr_en),
.number_out(VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2_number),
.read_add(VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2_read_add),
.data_out(VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI1X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X1;
wire PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X1_wr_en;
wire [5:0] VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1_number;
wire [8:0] VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1_read_add;
wire [13:0] VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1;
VMProjections  VMPROJ_F3F4_F2D5PHI2X1(
.data_in(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X1),
.enable(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X1_wr_en),
.number_out(VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1_number),
.read_add(VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1_read_add),
.data_out(VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1),
.start(PRD_F2D5_F3F4_start),
.done(VMPROJ_F3F4_F2D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI2X1n3;
wire VMRD_F2D5_VMS_F2D5PHI2X1n3_wr_en;
wire [5:0] VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1_number;
wire [10:0] VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1_read_add;
wire [18:0] VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1;
VMStubs #("Match") VMS_F2D5PHI2X1n3(
.data_in(VMRD_F2D5_VMS_F2D5PHI2X1n3),
.enable(VMRD_F2D5_VMS_F2D5PHI2X1n3_wr_en),
.number_out(VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1_number),
.read_add(VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1_read_add),
.data_out(VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X2;
wire PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X2_wr_en;
wire [5:0] VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2_number;
wire [8:0] VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2_read_add;
wire [13:0] VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2;
VMProjections  VMPROJ_F3F4_F2D5PHI2X2(
.data_in(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X2),
.enable(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X2_wr_en),
.number_out(VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2_number),
.read_add(VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2_read_add),
.data_out(VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2),
.start(PRD_F2D5_F3F4_start),
.done(VMPROJ_F3F4_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI2X2n5;
wire VMRD_F2D5_VMS_F2D5PHI2X2n5_wr_en;
wire [5:0] VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2_number;
wire [10:0] VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2_read_add;
wire [18:0] VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2;
VMStubs #("Match") VMS_F2D5PHI2X2n5(
.data_in(VMRD_F2D5_VMS_F2D5PHI2X2n5),
.enable(VMRD_F2D5_VMS_F2D5PHI2X2n5_wr_en),
.number_out(VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2_number),
.read_add(VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2_read_add),
.data_out(VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X1;
wire PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X1_wr_en;
wire [5:0] VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1_number;
wire [8:0] VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1_read_add;
wire [13:0] VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1;
VMProjections  VMPROJ_F3F4_F2D5PHI3X1(
.data_in(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X1),
.enable(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X1_wr_en),
.number_out(VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1_number),
.read_add(VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1_read_add),
.data_out(VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1),
.start(PRD_F2D5_F3F4_start),
.done(VMPROJ_F3F4_F2D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI3X1n3;
wire VMRD_F2D5_VMS_F2D5PHI3X1n3_wr_en;
wire [5:0] VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1_number;
wire [10:0] VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1_read_add;
wire [18:0] VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1;
VMStubs #("Match") VMS_F2D5PHI3X1n3(
.data_in(VMRD_F2D5_VMS_F2D5PHI3X1n3),
.enable(VMRD_F2D5_VMS_F2D5PHI3X1n3_wr_en),
.number_out(VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1_number),
.read_add(VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1_read_add),
.data_out(VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X2;
wire PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X2_wr_en;
wire [5:0] VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2_number;
wire [8:0] VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2_read_add;
wire [13:0] VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2;
VMProjections  VMPROJ_F3F4_F2D5PHI3X2(
.data_in(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X2),
.enable(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X2_wr_en),
.number_out(VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2_number),
.read_add(VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2_read_add),
.data_out(VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2),
.start(PRD_F2D5_F3F4_start),
.done(VMPROJ_F3F4_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F2D5_VMS_F2D5PHI3X2n5;
wire VMRD_F2D5_VMS_F2D5PHI3X2n5_wr_en;
wire [5:0] VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2_number;
wire [10:0] VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2_read_add;
wire [18:0] VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2;
VMStubs #("Match") VMS_F2D5PHI3X2n5(
.data_in(VMRD_F2D5_VMS_F2D5PHI3X2n5),
.enable(VMRD_F2D5_VMS_F2D5PHI3X2n5_wr_en),
.number_out(VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2_number),
.read_add(VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2_read_add),
.data_out(VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2),
.start(VMRD_F2D5_start),
.done(VMS_F2D5PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X1;
wire PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X1_wr_en;
wire [5:0] VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1_number;
wire [8:0] VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1_read_add;
wire [13:0] VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1;
VMProjections  VMPROJ_F3F4_F5D5PHI1X1(
.data_in(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X1),
.enable(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X1_wr_en),
.number_out(VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1_number),
.read_add(VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1_read_add),
.data_out(VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1),
.start(PRD_F5D5_F3F4_start),
.done(VMPROJ_F3F4_F5D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI1X1n2;
wire VMRD_F5D5_VMS_F5D5PHI1X1n2_wr_en;
wire [5:0] VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1_number;
wire [10:0] VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1_read_add;
wire [18:0] VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1;
VMStubs #("Match") VMS_F5D5PHI1X1n2(
.data_in(VMRD_F5D5_VMS_F5D5PHI1X1n2),
.enable(VMRD_F5D5_VMS_F5D5PHI1X1n2_wr_en),
.number_out(VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1_number),
.read_add(VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1_read_add),
.data_out(VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X2;
wire PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X2_wr_en;
wire [5:0] VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2_number;
wire [8:0] VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2_read_add;
wire [13:0] VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2;
VMProjections  VMPROJ_F3F4_F5D5PHI1X2(
.data_in(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X2),
.enable(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X2_wr_en),
.number_out(VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2_number),
.read_add(VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2_read_add),
.data_out(VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2),
.start(PRD_F5D5_F3F4_start),
.done(VMPROJ_F3F4_F5D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI1X2n2;
wire VMRD_F5D5_VMS_F5D5PHI1X2n2_wr_en;
wire [5:0] VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2_number;
wire [10:0] VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2_read_add;
wire [18:0] VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2;
VMStubs #("Match") VMS_F5D5PHI1X2n2(
.data_in(VMRD_F5D5_VMS_F5D5PHI1X2n2),
.enable(VMRD_F5D5_VMS_F5D5PHI1X2n2_wr_en),
.number_out(VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2_number),
.read_add(VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2_read_add),
.data_out(VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X1;
wire PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X1_wr_en;
wire [5:0] VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1_number;
wire [8:0] VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1_read_add;
wire [13:0] VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1;
VMProjections  VMPROJ_F3F4_F5D5PHI2X1(
.data_in(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X1),
.enable(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X1_wr_en),
.number_out(VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1_number),
.read_add(VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1_read_add),
.data_out(VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1),
.start(PRD_F5D5_F3F4_start),
.done(VMPROJ_F3F4_F5D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI2X1n2;
wire VMRD_F5D5_VMS_F5D5PHI2X1n2_wr_en;
wire [5:0] VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1_number;
wire [10:0] VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1_read_add;
wire [18:0] VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1;
VMStubs #("Match") VMS_F5D5PHI2X1n2(
.data_in(VMRD_F5D5_VMS_F5D5PHI2X1n2),
.enable(VMRD_F5D5_VMS_F5D5PHI2X1n2_wr_en),
.number_out(VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1_number),
.read_add(VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1_read_add),
.data_out(VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X2;
wire PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X2_wr_en;
wire [5:0] VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2_number;
wire [8:0] VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2_read_add;
wire [13:0] VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2;
VMProjections  VMPROJ_F3F4_F5D5PHI2X2(
.data_in(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X2),
.enable(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X2_wr_en),
.number_out(VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2_number),
.read_add(VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2_read_add),
.data_out(VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2),
.start(PRD_F5D5_F3F4_start),
.done(VMPROJ_F3F4_F5D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI2X2n2;
wire VMRD_F5D5_VMS_F5D5PHI2X2n2_wr_en;
wire [5:0] VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2_number;
wire [10:0] VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2_read_add;
wire [18:0] VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2;
VMStubs #("Match") VMS_F5D5PHI2X2n2(
.data_in(VMRD_F5D5_VMS_F5D5PHI2X2n2),
.enable(VMRD_F5D5_VMS_F5D5PHI2X2n2_wr_en),
.number_out(VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2_number),
.read_add(VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2_read_add),
.data_out(VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X1;
wire PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X1_wr_en;
wire [5:0] VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1_number;
wire [8:0] VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1_read_add;
wire [13:0] VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1;
VMProjections  VMPROJ_F3F4_F5D5PHI3X1(
.data_in(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X1),
.enable(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X1_wr_en),
.number_out(VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1_number),
.read_add(VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1_read_add),
.data_out(VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1),
.start(PRD_F5D5_F3F4_start),
.done(VMPROJ_F3F4_F5D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI3X1n2;
wire VMRD_F5D5_VMS_F5D5PHI3X1n2_wr_en;
wire [5:0] VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1_number;
wire [10:0] VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1_read_add;
wire [18:0] VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1;
VMStubs #("Match") VMS_F5D5PHI3X1n2(
.data_in(VMRD_F5D5_VMS_F5D5PHI3X1n2),
.enable(VMRD_F5D5_VMS_F5D5PHI3X1n2_wr_en),
.number_out(VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1_number),
.read_add(VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1_read_add),
.data_out(VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X2;
wire PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X2_wr_en;
wire [5:0] VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2_number;
wire [8:0] VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2_read_add;
wire [13:0] VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2;
VMProjections  VMPROJ_F3F4_F5D5PHI3X2(
.data_in(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X2),
.enable(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X2_wr_en),
.number_out(VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2_number),
.read_add(VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2_read_add),
.data_out(VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2),
.start(PRD_F5D5_F3F4_start),
.done(VMPROJ_F3F4_F5D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI3X2n2;
wire VMRD_F5D5_VMS_F5D5PHI3X2n2_wr_en;
wire [5:0] VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2_number;
wire [10:0] VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2_read_add;
wire [18:0] VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2;
VMStubs #("Match") VMS_F5D5PHI3X2n2(
.data_in(VMRD_F5D5_VMS_F5D5PHI3X2n2),
.enable(VMRD_F5D5_VMS_F5D5PHI3X2n2_wr_en),
.number_out(VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2_number),
.read_add(VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2_read_add),
.data_out(VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X1;
wire PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X1_wr_en;
wire [5:0] VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1_number;
wire [8:0] VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1_read_add;
wire [13:0] VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1;
VMProjections  VMPROJ_F3F4_F5D5PHI4X1(
.data_in(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X1),
.enable(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X1_wr_en),
.number_out(VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1_number),
.read_add(VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1_read_add),
.data_out(VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1),
.start(PRD_F5D5_F3F4_start),
.done(VMPROJ_F3F4_F5D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI4X1n2;
wire VMRD_F5D5_VMS_F5D5PHI4X1n2_wr_en;
wire [5:0] VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1_number;
wire [10:0] VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1_read_add;
wire [18:0] VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1;
VMStubs #("Match") VMS_F5D5PHI4X1n2(
.data_in(VMRD_F5D5_VMS_F5D5PHI4X1n2),
.enable(VMRD_F5D5_VMS_F5D5PHI4X1n2_wr_en),
.number_out(VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1_number),
.read_add(VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1_read_add),
.data_out(VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X2;
wire PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X2_wr_en;
wire [5:0] VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2_number;
wire [8:0] VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2_read_add;
wire [13:0] VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2;
VMProjections  VMPROJ_F3F4_F5D5PHI4X2(
.data_in(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X2),
.enable(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X2_wr_en),
.number_out(VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2_number),
.read_add(VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2_read_add),
.data_out(VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2),
.start(PRD_F5D5_F3F4_start),
.done(VMPROJ_F3F4_F5D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMRD_F5D5_VMS_F5D5PHI4X2n2;
wire VMRD_F5D5_VMS_F5D5PHI4X2n2_wr_en;
wire [5:0] VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2_number;
wire [10:0] VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2_read_add;
wire [18:0] VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2;
VMStubs #("Match") VMS_F5D5PHI4X2n2(
.data_in(VMRD_F5D5_VMS_F5D5PHI4X2n2),
.enable(VMRD_F5D5_VMS_F5D5PHI4X2n2_wr_en),
.number_out(VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2_number),
.read_add(VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2_read_add),
.data_out(VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2),
.start(VMRD_F5D5_start),
.done(VMS_F5D5PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F3D5PHI1X1_CM_F1F2_F3D5PHI1X1;
wire ME_F1F2_F3D5PHI1X1_CM_F1F2_F3D5PHI1X1_wr_en;
wire [5:0] CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5_number;
wire [8:0] CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5_read_add;
wire [11:0] CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5;
CandidateMatch  CM_F1F2_F3D5PHI1X1(
.data_in(ME_F1F2_F3D5PHI1X1_CM_F1F2_F3D5PHI1X1),
.enable(ME_F1F2_F3D5PHI1X1_CM_F1F2_F3D5PHI1X1_wr_en),
.number_out(CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5_number),
.read_add(CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5_read_add),
.data_out(CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5),
.start(ME_F1F2_F3D5PHI1X1_start),
.done(CM_F1F2_F3D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F3D5PHI1X2_CM_F1F2_F3D5PHI1X2;
wire ME_F1F2_F3D5PHI1X2_CM_F1F2_F3D5PHI1X2_wr_en;
wire [5:0] CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5_number;
wire [8:0] CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5_read_add;
wire [11:0] CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5;
CandidateMatch  CM_F1F2_F3D5PHI1X2(
.data_in(ME_F1F2_F3D5PHI1X2_CM_F1F2_F3D5PHI1X2),
.enable(ME_F1F2_F3D5PHI1X2_CM_F1F2_F3D5PHI1X2_wr_en),
.number_out(CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5_number),
.read_add(CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5_read_add),
.data_out(CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5),
.start(ME_F1F2_F3D5PHI1X2_start),
.done(CM_F1F2_F3D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F3D5PHI2X1_CM_F1F2_F3D5PHI2X1;
wire ME_F1F2_F3D5PHI2X1_CM_F1F2_F3D5PHI2X1_wr_en;
wire [5:0] CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5_number;
wire [8:0] CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5_read_add;
wire [11:0] CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5;
CandidateMatch  CM_F1F2_F3D5PHI2X1(
.data_in(ME_F1F2_F3D5PHI2X1_CM_F1F2_F3D5PHI2X1),
.enable(ME_F1F2_F3D5PHI2X1_CM_F1F2_F3D5PHI2X1_wr_en),
.number_out(CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5_number),
.read_add(CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5_read_add),
.data_out(CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5),
.start(ME_F1F2_F3D5PHI2X1_start),
.done(CM_F1F2_F3D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F3D5PHI2X2_CM_F1F2_F3D5PHI2X2;
wire ME_F1F2_F3D5PHI2X2_CM_F1F2_F3D5PHI2X2_wr_en;
wire [5:0] CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5_number;
wire [8:0] CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5_read_add;
wire [11:0] CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5;
CandidateMatch  CM_F1F2_F3D5PHI2X2(
.data_in(ME_F1F2_F3D5PHI2X2_CM_F1F2_F3D5PHI2X2),
.enable(ME_F1F2_F3D5PHI2X2_CM_F1F2_F3D5PHI2X2_wr_en),
.number_out(CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5_number),
.read_add(CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5_read_add),
.data_out(CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5),
.start(ME_F1F2_F3D5PHI2X2_start),
.done(CM_F1F2_F3D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F3D5PHI3X1_CM_F1F2_F3D5PHI3X1;
wire ME_F1F2_F3D5PHI3X1_CM_F1F2_F3D5PHI3X1_wr_en;
wire [5:0] CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5_number;
wire [8:0] CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5_read_add;
wire [11:0] CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5;
CandidateMatch  CM_F1F2_F3D5PHI3X1(
.data_in(ME_F1F2_F3D5PHI3X1_CM_F1F2_F3D5PHI3X1),
.enable(ME_F1F2_F3D5PHI3X1_CM_F1F2_F3D5PHI3X1_wr_en),
.number_out(CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5_number),
.read_add(CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5_read_add),
.data_out(CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5),
.start(ME_F1F2_F3D5PHI3X1_start),
.done(CM_F1F2_F3D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F3D5PHI3X2_CM_F1F2_F3D5PHI3X2;
wire ME_F1F2_F3D5PHI3X2_CM_F1F2_F3D5PHI3X2_wr_en;
wire [5:0] CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5_number;
wire [8:0] CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5_read_add;
wire [11:0] CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5;
CandidateMatch  CM_F1F2_F3D5PHI3X2(
.data_in(ME_F1F2_F3D5PHI3X2_CM_F1F2_F3D5PHI3X2),
.enable(ME_F1F2_F3D5PHI3X2_CM_F1F2_F3D5PHI3X2_wr_en),
.number_out(CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5_number),
.read_add(CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5_read_add),
.data_out(CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5),
.start(ME_F1F2_F3D5PHI3X2_start),
.done(CM_F1F2_F3D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F3D5PHI4X1_CM_F1F2_F3D5PHI4X1;
wire ME_F1F2_F3D5PHI4X1_CM_F1F2_F3D5PHI4X1_wr_en;
wire [5:0] CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5_number;
wire [8:0] CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5_read_add;
wire [11:0] CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5;
CandidateMatch  CM_F1F2_F3D5PHI4X1(
.data_in(ME_F1F2_F3D5PHI4X1_CM_F1F2_F3D5PHI4X1),
.enable(ME_F1F2_F3D5PHI4X1_CM_F1F2_F3D5PHI4X1_wr_en),
.number_out(CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5_number),
.read_add(CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5_read_add),
.data_out(CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5),
.start(ME_F1F2_F3D5PHI4X1_start),
.done(CM_F1F2_F3D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F3D5PHI4X2_CM_F1F2_F3D5PHI4X2;
wire ME_F1F2_F3D5PHI4X2_CM_F1F2_F3D5PHI4X2_wr_en;
wire [5:0] CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5_number;
wire [8:0] CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5_read_add;
wire [11:0] CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5;
CandidateMatch  CM_F1F2_F3D5PHI4X2(
.data_in(ME_F1F2_F3D5PHI4X2_CM_F1F2_F3D5PHI4X2),
.enable(ME_F1F2_F3D5PHI4X2_CM_F1F2_F3D5PHI4X2_wr_en),
.number_out(CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5_number),
.read_add(CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5_read_add),
.data_out(CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5),
.start(ME_F1F2_F3D5PHI4X2_start),
.done(CM_F1F2_F3D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PRD_F3D5_F1F2_AP_F1F2_F3D5;
wire PRD_F3D5_F1F2_AP_F1F2_F3D5_wr_en;
wire [8:0] AP_F1F2_F3D5_MC_F1F2_F3D5_read_add;
wire [55:0] AP_F1F2_F3D5_MC_F1F2_F3D5;
AllProj #(1'b0,1'b1) AP_F1F2_F3D5(
.data_in(PRD_F3D5_F1F2_AP_F1F2_F3D5),
.enable(PRD_F3D5_F1F2_AP_F1F2_F3D5_wr_en),
.read_add(AP_F1F2_F3D5_MC_F1F2_F3D5_read_add),
.data_out(AP_F1F2_F3D5_MC_F1F2_F3D5),
.start(PRD_F3D5_F1F2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F3D5_AS_F3D5n2;
wire VMRD_F3D5_AS_F3D5n2_wr_en;
wire [10:0] AS_F3D5n2_MC_F1F2_F3D5_read_add;
wire [35:0] AS_F3D5n2_MC_F1F2_F3D5;
AllStubs  AS_F3D5n2(
.data_in(VMRD_F3D5_AS_F3D5n2),
.enable(VMRD_F3D5_AS_F3D5n2_wr_en),
.read_add_MC(AS_F3D5n2_MC_F1F2_F3D5_read_add),
.data_out_MC(AS_F3D5n2_MC_F1F2_F3D5),
.start(VMRD_F3D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F4D5PHI1X1_CM_F1F2_F4D5PHI1X1;
wire ME_F1F2_F4D5PHI1X1_CM_F1F2_F4D5PHI1X1_wr_en;
wire [5:0] CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5_number;
wire [8:0] CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5_read_add;
wire [11:0] CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5;
CandidateMatch  CM_F1F2_F4D5PHI1X1(
.data_in(ME_F1F2_F4D5PHI1X1_CM_F1F2_F4D5PHI1X1),
.enable(ME_F1F2_F4D5PHI1X1_CM_F1F2_F4D5PHI1X1_wr_en),
.number_out(CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5_number),
.read_add(CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5_read_add),
.data_out(CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5),
.start(ME_F1F2_F4D5PHI1X1_start),
.done(CM_F1F2_F4D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F4D5PHI1X2_CM_F1F2_F4D5PHI1X2;
wire ME_F1F2_F4D5PHI1X2_CM_F1F2_F4D5PHI1X2_wr_en;
wire [5:0] CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5_number;
wire [8:0] CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5_read_add;
wire [11:0] CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5;
CandidateMatch  CM_F1F2_F4D5PHI1X2(
.data_in(ME_F1F2_F4D5PHI1X2_CM_F1F2_F4D5PHI1X2),
.enable(ME_F1F2_F4D5PHI1X2_CM_F1F2_F4D5PHI1X2_wr_en),
.number_out(CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5_number),
.read_add(CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5_read_add),
.data_out(CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5),
.start(ME_F1F2_F4D5PHI1X2_start),
.done(CM_F1F2_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F4D5PHI2X1_CM_F1F2_F4D5PHI2X1;
wire ME_F1F2_F4D5PHI2X1_CM_F1F2_F4D5PHI2X1_wr_en;
wire [5:0] CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5_number;
wire [8:0] CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5_read_add;
wire [11:0] CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5;
CandidateMatch  CM_F1F2_F4D5PHI2X1(
.data_in(ME_F1F2_F4D5PHI2X1_CM_F1F2_F4D5PHI2X1),
.enable(ME_F1F2_F4D5PHI2X1_CM_F1F2_F4D5PHI2X1_wr_en),
.number_out(CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5_number),
.read_add(CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5_read_add),
.data_out(CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5),
.start(ME_F1F2_F4D5PHI2X1_start),
.done(CM_F1F2_F4D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F4D5PHI2X2_CM_F1F2_F4D5PHI2X2;
wire ME_F1F2_F4D5PHI2X2_CM_F1F2_F4D5PHI2X2_wr_en;
wire [5:0] CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5_number;
wire [8:0] CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5_read_add;
wire [11:0] CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5;
CandidateMatch  CM_F1F2_F4D5PHI2X2(
.data_in(ME_F1F2_F4D5PHI2X2_CM_F1F2_F4D5PHI2X2),
.enable(ME_F1F2_F4D5PHI2X2_CM_F1F2_F4D5PHI2X2_wr_en),
.number_out(CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5_number),
.read_add(CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5_read_add),
.data_out(CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5),
.start(ME_F1F2_F4D5PHI2X2_start),
.done(CM_F1F2_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F4D5PHI3X1_CM_F1F2_F4D5PHI3X1;
wire ME_F1F2_F4D5PHI3X1_CM_F1F2_F4D5PHI3X1_wr_en;
wire [5:0] CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5_number;
wire [8:0] CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5_read_add;
wire [11:0] CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5;
CandidateMatch  CM_F1F2_F4D5PHI3X1(
.data_in(ME_F1F2_F4D5PHI3X1_CM_F1F2_F4D5PHI3X1),
.enable(ME_F1F2_F4D5PHI3X1_CM_F1F2_F4D5PHI3X1_wr_en),
.number_out(CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5_number),
.read_add(CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5_read_add),
.data_out(CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5),
.start(ME_F1F2_F4D5PHI3X1_start),
.done(CM_F1F2_F4D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F4D5PHI3X2_CM_F1F2_F4D5PHI3X2;
wire ME_F1F2_F4D5PHI3X2_CM_F1F2_F4D5PHI3X2_wr_en;
wire [5:0] CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5_number;
wire [8:0] CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5_read_add;
wire [11:0] CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5;
CandidateMatch  CM_F1F2_F4D5PHI3X2(
.data_in(ME_F1F2_F4D5PHI3X2_CM_F1F2_F4D5PHI3X2),
.enable(ME_F1F2_F4D5PHI3X2_CM_F1F2_F4D5PHI3X2_wr_en),
.number_out(CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5_number),
.read_add(CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5_read_add),
.data_out(CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5),
.start(ME_F1F2_F4D5PHI3X2_start),
.done(CM_F1F2_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PRD_F4D5_F1F2_AP_F1F2_F4D5;
wire PRD_F4D5_F1F2_AP_F1F2_F4D5_wr_en;
wire [8:0] AP_F1F2_F4D5_MC_F1F2_F4D5_read_add;
wire [55:0] AP_F1F2_F4D5_MC_F1F2_F4D5;
AllProj #(1'b0,1'b1) AP_F1F2_F4D5(
.data_in(PRD_F4D5_F1F2_AP_F1F2_F4D5),
.enable(PRD_F4D5_F1F2_AP_F1F2_F4D5_wr_en),
.read_add(AP_F1F2_F4D5_MC_F1F2_F4D5_read_add),
.data_out(AP_F1F2_F4D5_MC_F1F2_F4D5),
.start(PRD_F4D5_F1F2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F4D5_AS_F4D5n2;
wire VMRD_F4D5_AS_F4D5n2_wr_en;
wire [10:0] AS_F4D5n2_MC_F1F2_F4D5_read_add;
wire [35:0] AS_F4D5n2_MC_F1F2_F4D5;
AllStubs  AS_F4D5n2(
.data_in(VMRD_F4D5_AS_F4D5n2),
.enable(VMRD_F4D5_AS_F4D5n2_wr_en),
.read_add_MC(AS_F4D5n2_MC_F1F2_F4D5_read_add),
.data_out_MC(AS_F4D5n2_MC_F1F2_F4D5),
.start(VMRD_F4D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F5D5PHI1X1_CM_F1F2_F5D5PHI1X1;
wire ME_F1F2_F5D5PHI1X1_CM_F1F2_F5D5PHI1X1_wr_en;
wire [5:0] CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5_number;
wire [8:0] CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5_read_add;
wire [11:0] CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5;
CandidateMatch  CM_F1F2_F5D5PHI1X1(
.data_in(ME_F1F2_F5D5PHI1X1_CM_F1F2_F5D5PHI1X1),
.enable(ME_F1F2_F5D5PHI1X1_CM_F1F2_F5D5PHI1X1_wr_en),
.number_out(CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5_number),
.read_add(CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5_read_add),
.data_out(CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5),
.start(ME_F1F2_F5D5PHI1X1_start),
.done(CM_F1F2_F5D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F5D5PHI1X2_CM_F1F2_F5D5PHI1X2;
wire ME_F1F2_F5D5PHI1X2_CM_F1F2_F5D5PHI1X2_wr_en;
wire [5:0] CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5_number;
wire [8:0] CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5_read_add;
wire [11:0] CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5;
CandidateMatch  CM_F1F2_F5D5PHI1X2(
.data_in(ME_F1F2_F5D5PHI1X2_CM_F1F2_F5D5PHI1X2),
.enable(ME_F1F2_F5D5PHI1X2_CM_F1F2_F5D5PHI1X2_wr_en),
.number_out(CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5_number),
.read_add(CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5_read_add),
.data_out(CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5),
.start(ME_F1F2_F5D5PHI1X2_start),
.done(CM_F1F2_F5D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F5D5PHI2X1_CM_F1F2_F5D5PHI2X1;
wire ME_F1F2_F5D5PHI2X1_CM_F1F2_F5D5PHI2X1_wr_en;
wire [5:0] CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5_number;
wire [8:0] CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5_read_add;
wire [11:0] CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5;
CandidateMatch  CM_F1F2_F5D5PHI2X1(
.data_in(ME_F1F2_F5D5PHI2X1_CM_F1F2_F5D5PHI2X1),
.enable(ME_F1F2_F5D5PHI2X1_CM_F1F2_F5D5PHI2X1_wr_en),
.number_out(CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5_number),
.read_add(CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5_read_add),
.data_out(CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5),
.start(ME_F1F2_F5D5PHI2X1_start),
.done(CM_F1F2_F5D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F5D5PHI2X2_CM_F1F2_F5D5PHI2X2;
wire ME_F1F2_F5D5PHI2X2_CM_F1F2_F5D5PHI2X2_wr_en;
wire [5:0] CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5_number;
wire [8:0] CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5_read_add;
wire [11:0] CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5;
CandidateMatch  CM_F1F2_F5D5PHI2X2(
.data_in(ME_F1F2_F5D5PHI2X2_CM_F1F2_F5D5PHI2X2),
.enable(ME_F1F2_F5D5PHI2X2_CM_F1F2_F5D5PHI2X2_wr_en),
.number_out(CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5_number),
.read_add(CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5_read_add),
.data_out(CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5),
.start(ME_F1F2_F5D5PHI2X2_start),
.done(CM_F1F2_F5D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F5D5PHI3X1_CM_F1F2_F5D5PHI3X1;
wire ME_F1F2_F5D5PHI3X1_CM_F1F2_F5D5PHI3X1_wr_en;
wire [5:0] CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5_number;
wire [8:0] CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5_read_add;
wire [11:0] CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5;
CandidateMatch  CM_F1F2_F5D5PHI3X1(
.data_in(ME_F1F2_F5D5PHI3X1_CM_F1F2_F5D5PHI3X1),
.enable(ME_F1F2_F5D5PHI3X1_CM_F1F2_F5D5PHI3X1_wr_en),
.number_out(CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5_number),
.read_add(CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5_read_add),
.data_out(CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5),
.start(ME_F1F2_F5D5PHI3X1_start),
.done(CM_F1F2_F5D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F5D5PHI3X2_CM_F1F2_F5D5PHI3X2;
wire ME_F1F2_F5D5PHI3X2_CM_F1F2_F5D5PHI3X2_wr_en;
wire [5:0] CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5_number;
wire [8:0] CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5_read_add;
wire [11:0] CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5;
CandidateMatch  CM_F1F2_F5D5PHI3X2(
.data_in(ME_F1F2_F5D5PHI3X2_CM_F1F2_F5D5PHI3X2),
.enable(ME_F1F2_F5D5PHI3X2_CM_F1F2_F5D5PHI3X2_wr_en),
.number_out(CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5_number),
.read_add(CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5_read_add),
.data_out(CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5),
.start(ME_F1F2_F5D5PHI3X2_start),
.done(CM_F1F2_F5D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F5D5PHI4X1_CM_F1F2_F5D5PHI4X1;
wire ME_F1F2_F5D5PHI4X1_CM_F1F2_F5D5PHI4X1_wr_en;
wire [5:0] CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5_number;
wire [8:0] CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5_read_add;
wire [11:0] CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5;
CandidateMatch  CM_F1F2_F5D5PHI4X1(
.data_in(ME_F1F2_F5D5PHI4X1_CM_F1F2_F5D5PHI4X1),
.enable(ME_F1F2_F5D5PHI4X1_CM_F1F2_F5D5PHI4X1_wr_en),
.number_out(CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5_number),
.read_add(CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5_read_add),
.data_out(CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5),
.start(ME_F1F2_F5D5PHI4X1_start),
.done(CM_F1F2_F5D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F1F2_F5D5PHI4X2_CM_F1F2_F5D5PHI4X2;
wire ME_F1F2_F5D5PHI4X2_CM_F1F2_F5D5PHI4X2_wr_en;
wire [5:0] CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5_number;
wire [8:0] CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5_read_add;
wire [11:0] CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5;
CandidateMatch  CM_F1F2_F5D5PHI4X2(
.data_in(ME_F1F2_F5D5PHI4X2_CM_F1F2_F5D5PHI4X2),
.enable(ME_F1F2_F5D5PHI4X2_CM_F1F2_F5D5PHI4X2_wr_en),
.number_out(CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5_number),
.read_add(CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5_read_add),
.data_out(CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5),
.start(ME_F1F2_F5D5PHI4X2_start),
.done(CM_F1F2_F5D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PRD_F5D5_F1F2_AP_F1F2_F5D5;
wire PRD_F5D5_F1F2_AP_F1F2_F5D5_wr_en;
wire [8:0] AP_F1F2_F5D5_MC_F1F2_F5D5_read_add;
wire [55:0] AP_F1F2_F5D5_MC_F1F2_F5D5;
AllProj #(1'b0,1'b1) AP_F1F2_F5D5(
.data_in(PRD_F5D5_F1F2_AP_F1F2_F5D5),
.enable(PRD_F5D5_F1F2_AP_F1F2_F5D5_wr_en),
.read_add(AP_F1F2_F5D5_MC_F1F2_F5D5_read_add),
.data_out(AP_F1F2_F5D5_MC_F1F2_F5D5),
.start(PRD_F5D5_F1F2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F5D5_AS_F5D5n1;
wire VMRD_F5D5_AS_F5D5n1_wr_en;
wire [10:0] AS_F5D5n1_MC_F1F2_F5D5_read_add;
wire [35:0] AS_F5D5n1_MC_F1F2_F5D5;
AllStubs  AS_F5D5n1(
.data_in(VMRD_F5D5_AS_F5D5n1),
.enable(VMRD_F5D5_AS_F5D5n1_wr_en),
.read_add_MC(AS_F5D5n1_MC_F1F2_F5D5_read_add),
.data_out_MC(AS_F5D5n1_MC_F1F2_F5D5),
.start(VMRD_F5D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F1D5PHI1X1_CM_F3F4_F1D5PHI1X1;
wire ME_F3F4_F1D5PHI1X1_CM_F3F4_F1D5PHI1X1_wr_en;
wire [5:0] CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5_number;
wire [8:0] CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5_read_add;
wire [11:0] CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5;
CandidateMatch  CM_F3F4_F1D5PHI1X1(
.data_in(ME_F3F4_F1D5PHI1X1_CM_F3F4_F1D5PHI1X1),
.enable(ME_F3F4_F1D5PHI1X1_CM_F3F4_F1D5PHI1X1_wr_en),
.number_out(CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5_number),
.read_add(CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5_read_add),
.data_out(CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5),
.start(ME_F3F4_F1D5PHI1X1_start),
.done(CM_F3F4_F1D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F1D5PHI1X2_CM_F3F4_F1D5PHI1X2;
wire ME_F3F4_F1D5PHI1X2_CM_F3F4_F1D5PHI1X2_wr_en;
wire [5:0] CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5_number;
wire [8:0] CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5_read_add;
wire [11:0] CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5;
CandidateMatch  CM_F3F4_F1D5PHI1X2(
.data_in(ME_F3F4_F1D5PHI1X2_CM_F3F4_F1D5PHI1X2),
.enable(ME_F3F4_F1D5PHI1X2_CM_F3F4_F1D5PHI1X2_wr_en),
.number_out(CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5_number),
.read_add(CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5_read_add),
.data_out(CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5),
.start(ME_F3F4_F1D5PHI1X2_start),
.done(CM_F3F4_F1D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F1D5PHI2X1_CM_F3F4_F1D5PHI2X1;
wire ME_F3F4_F1D5PHI2X1_CM_F3F4_F1D5PHI2X1_wr_en;
wire [5:0] CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5_number;
wire [8:0] CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5_read_add;
wire [11:0] CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5;
CandidateMatch  CM_F3F4_F1D5PHI2X1(
.data_in(ME_F3F4_F1D5PHI2X1_CM_F3F4_F1D5PHI2X1),
.enable(ME_F3F4_F1D5PHI2X1_CM_F3F4_F1D5PHI2X1_wr_en),
.number_out(CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5_number),
.read_add(CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5_read_add),
.data_out(CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5),
.start(ME_F3F4_F1D5PHI2X1_start),
.done(CM_F3F4_F1D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F1D5PHI2X2_CM_F3F4_F1D5PHI2X2;
wire ME_F3F4_F1D5PHI2X2_CM_F3F4_F1D5PHI2X2_wr_en;
wire [5:0] CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5_number;
wire [8:0] CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5_read_add;
wire [11:0] CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5;
CandidateMatch  CM_F3F4_F1D5PHI2X2(
.data_in(ME_F3F4_F1D5PHI2X2_CM_F3F4_F1D5PHI2X2),
.enable(ME_F3F4_F1D5PHI2X2_CM_F3F4_F1D5PHI2X2_wr_en),
.number_out(CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5_number),
.read_add(CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5_read_add),
.data_out(CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5),
.start(ME_F3F4_F1D5PHI2X2_start),
.done(CM_F3F4_F1D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F1D5PHI3X1_CM_F3F4_F1D5PHI3X1;
wire ME_F3F4_F1D5PHI3X1_CM_F3F4_F1D5PHI3X1_wr_en;
wire [5:0] CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5_number;
wire [8:0] CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5_read_add;
wire [11:0] CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5;
CandidateMatch  CM_F3F4_F1D5PHI3X1(
.data_in(ME_F3F4_F1D5PHI3X1_CM_F3F4_F1D5PHI3X1),
.enable(ME_F3F4_F1D5PHI3X1_CM_F3F4_F1D5PHI3X1_wr_en),
.number_out(CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5_number),
.read_add(CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5_read_add),
.data_out(CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5),
.start(ME_F3F4_F1D5PHI3X1_start),
.done(CM_F3F4_F1D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F1D5PHI3X2_CM_F3F4_F1D5PHI3X2;
wire ME_F3F4_F1D5PHI3X2_CM_F3F4_F1D5PHI3X2_wr_en;
wire [5:0] CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5_number;
wire [8:0] CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5_read_add;
wire [11:0] CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5;
CandidateMatch  CM_F3F4_F1D5PHI3X2(
.data_in(ME_F3F4_F1D5PHI3X2_CM_F3F4_F1D5PHI3X2),
.enable(ME_F3F4_F1D5PHI3X2_CM_F3F4_F1D5PHI3X2_wr_en),
.number_out(CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5_number),
.read_add(CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5_read_add),
.data_out(CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5),
.start(ME_F3F4_F1D5PHI3X2_start),
.done(CM_F3F4_F1D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F1D5PHI4X1_CM_F3F4_F1D5PHI4X1;
wire ME_F3F4_F1D5PHI4X1_CM_F3F4_F1D5PHI4X1_wr_en;
wire [5:0] CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5_number;
wire [8:0] CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5_read_add;
wire [11:0] CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5;
CandidateMatch  CM_F3F4_F1D5PHI4X1(
.data_in(ME_F3F4_F1D5PHI4X1_CM_F3F4_F1D5PHI4X1),
.enable(ME_F3F4_F1D5PHI4X1_CM_F3F4_F1D5PHI4X1_wr_en),
.number_out(CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5_number),
.read_add(CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5_read_add),
.data_out(CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5),
.start(ME_F3F4_F1D5PHI4X1_start),
.done(CM_F3F4_F1D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F1D5PHI4X2_CM_F3F4_F1D5PHI4X2;
wire ME_F3F4_F1D5PHI4X2_CM_F3F4_F1D5PHI4X2_wr_en;
wire [5:0] CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5_number;
wire [8:0] CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5_read_add;
wire [11:0] CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5;
CandidateMatch  CM_F3F4_F1D5PHI4X2(
.data_in(ME_F3F4_F1D5PHI4X2_CM_F3F4_F1D5PHI4X2),
.enable(ME_F3F4_F1D5PHI4X2_CM_F3F4_F1D5PHI4X2_wr_en),
.number_out(CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5_number),
.read_add(CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5_read_add),
.data_out(CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5),
.start(ME_F3F4_F1D5PHI4X2_start),
.done(CM_F3F4_F1D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PRD_F1D5_F3F4_AP_F3F4_F1D5;
wire PRD_F1D5_F3F4_AP_F3F4_F1D5_wr_en;
wire [8:0] AP_F3F4_F1D5_MC_F3F4_F1D5_read_add;
wire [55:0] AP_F3F4_F1D5_MC_F3F4_F1D5;
AllProj #(1'b0,1'b1) AP_F3F4_F1D5(
.data_in(PRD_F1D5_F3F4_AP_F3F4_F1D5),
.enable(PRD_F1D5_F3F4_AP_F3F4_F1D5_wr_en),
.read_add(AP_F3F4_F1D5_MC_F3F4_F1D5_read_add),
.data_out(AP_F3F4_F1D5_MC_F3F4_F1D5),
.start(PRD_F1D5_F3F4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F1D5_AS_F1D5n2;
wire VMRD_F1D5_AS_F1D5n2_wr_en;
wire [10:0] AS_F1D5n2_MC_F3F4_F1D5_read_add;
wire [35:0] AS_F1D5n2_MC_F3F4_F1D5;
AllStubs  AS_F1D5n2(
.data_in(VMRD_F1D5_AS_F1D5n2),
.enable(VMRD_F1D5_AS_F1D5n2_wr_en),
.read_add_MC(AS_F1D5n2_MC_F3F4_F1D5_read_add),
.data_out_MC(AS_F1D5n2_MC_F3F4_F1D5),
.start(VMRD_F1D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F2D5PHI1X1_CM_F3F4_F2D5PHI1X1;
wire ME_F3F4_F2D5PHI1X1_CM_F3F4_F2D5PHI1X1_wr_en;
wire [5:0] CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5_number;
wire [8:0] CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5_read_add;
wire [11:0] CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5;
CandidateMatch  CM_F3F4_F2D5PHI1X1(
.data_in(ME_F3F4_F2D5PHI1X1_CM_F3F4_F2D5PHI1X1),
.enable(ME_F3F4_F2D5PHI1X1_CM_F3F4_F2D5PHI1X1_wr_en),
.number_out(CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5_number),
.read_add(CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5_read_add),
.data_out(CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5),
.start(ME_F3F4_F2D5PHI1X1_start),
.done(CM_F3F4_F2D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F2D5PHI1X2_CM_F3F4_F2D5PHI1X2;
wire ME_F3F4_F2D5PHI1X2_CM_F3F4_F2D5PHI1X2_wr_en;
wire [5:0] CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5_number;
wire [8:0] CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5_read_add;
wire [11:0] CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5;
CandidateMatch  CM_F3F4_F2D5PHI1X2(
.data_in(ME_F3F4_F2D5PHI1X2_CM_F3F4_F2D5PHI1X2),
.enable(ME_F3F4_F2D5PHI1X2_CM_F3F4_F2D5PHI1X2_wr_en),
.number_out(CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5_number),
.read_add(CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5_read_add),
.data_out(CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5),
.start(ME_F3F4_F2D5PHI1X2_start),
.done(CM_F3F4_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F2D5PHI2X1_CM_F3F4_F2D5PHI2X1;
wire ME_F3F4_F2D5PHI2X1_CM_F3F4_F2D5PHI2X1_wr_en;
wire [5:0] CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5_number;
wire [8:0] CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5_read_add;
wire [11:0] CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5;
CandidateMatch  CM_F3F4_F2D5PHI2X1(
.data_in(ME_F3F4_F2D5PHI2X1_CM_F3F4_F2D5PHI2X1),
.enable(ME_F3F4_F2D5PHI2X1_CM_F3F4_F2D5PHI2X1_wr_en),
.number_out(CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5_number),
.read_add(CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5_read_add),
.data_out(CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5),
.start(ME_F3F4_F2D5PHI2X1_start),
.done(CM_F3F4_F2D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F2D5PHI2X2_CM_F3F4_F2D5PHI2X2;
wire ME_F3F4_F2D5PHI2X2_CM_F3F4_F2D5PHI2X2_wr_en;
wire [5:0] CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5_number;
wire [8:0] CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5_read_add;
wire [11:0] CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5;
CandidateMatch  CM_F3F4_F2D5PHI2X2(
.data_in(ME_F3F4_F2D5PHI2X2_CM_F3F4_F2D5PHI2X2),
.enable(ME_F3F4_F2D5PHI2X2_CM_F3F4_F2D5PHI2X2_wr_en),
.number_out(CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5_number),
.read_add(CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5_read_add),
.data_out(CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5),
.start(ME_F3F4_F2D5PHI2X2_start),
.done(CM_F3F4_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F2D5PHI3X1_CM_F3F4_F2D5PHI3X1;
wire ME_F3F4_F2D5PHI3X1_CM_F3F4_F2D5PHI3X1_wr_en;
wire [5:0] CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5_number;
wire [8:0] CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5_read_add;
wire [11:0] CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5;
CandidateMatch  CM_F3F4_F2D5PHI3X1(
.data_in(ME_F3F4_F2D5PHI3X1_CM_F3F4_F2D5PHI3X1),
.enable(ME_F3F4_F2D5PHI3X1_CM_F3F4_F2D5PHI3X1_wr_en),
.number_out(CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5_number),
.read_add(CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5_read_add),
.data_out(CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5),
.start(ME_F3F4_F2D5PHI3X1_start),
.done(CM_F3F4_F2D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F2D5PHI3X2_CM_F3F4_F2D5PHI3X2;
wire ME_F3F4_F2D5PHI3X2_CM_F3F4_F2D5PHI3X2_wr_en;
wire [5:0] CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5_number;
wire [8:0] CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5_read_add;
wire [11:0] CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5;
CandidateMatch  CM_F3F4_F2D5PHI3X2(
.data_in(ME_F3F4_F2D5PHI3X2_CM_F3F4_F2D5PHI3X2),
.enable(ME_F3F4_F2D5PHI3X2_CM_F3F4_F2D5PHI3X2_wr_en),
.number_out(CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5_number),
.read_add(CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5_read_add),
.data_out(CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5),
.start(ME_F3F4_F2D5PHI3X2_start),
.done(CM_F3F4_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PRD_F2D5_F3F4_AP_F3F4_F2D5;
wire PRD_F2D5_F3F4_AP_F3F4_F2D5_wr_en;
wire [8:0] AP_F3F4_F2D5_MC_F3F4_F2D5_read_add;
wire [55:0] AP_F3F4_F2D5_MC_F3F4_F2D5;
AllProj #(1'b0,1'b1) AP_F3F4_F2D5(
.data_in(PRD_F2D5_F3F4_AP_F3F4_F2D5),
.enable(PRD_F2D5_F3F4_AP_F3F4_F2D5_wr_en),
.read_add(AP_F3F4_F2D5_MC_F3F4_F2D5_read_add),
.data_out(AP_F3F4_F2D5_MC_F3F4_F2D5),
.start(PRD_F2D5_F3F4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F2D5_AS_F2D5n2;
wire VMRD_F2D5_AS_F2D5n2_wr_en;
wire [10:0] AS_F2D5n2_MC_F3F4_F2D5_read_add;
wire [35:0] AS_F2D5n2_MC_F3F4_F2D5;
AllStubs  AS_F2D5n2(
.data_in(VMRD_F2D5_AS_F2D5n2),
.enable(VMRD_F2D5_AS_F2D5n2_wr_en),
.read_add_MC(AS_F2D5n2_MC_F3F4_F2D5_read_add),
.data_out_MC(AS_F2D5n2_MC_F3F4_F2D5),
.start(VMRD_F2D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F5D5PHI1X1_CM_F3F4_F5D5PHI1X1;
wire ME_F3F4_F5D5PHI1X1_CM_F3F4_F5D5PHI1X1_wr_en;
wire [5:0] CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5_number;
wire [8:0] CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5_read_add;
wire [11:0] CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5;
CandidateMatch  CM_F3F4_F5D5PHI1X1(
.data_in(ME_F3F4_F5D5PHI1X1_CM_F3F4_F5D5PHI1X1),
.enable(ME_F3F4_F5D5PHI1X1_CM_F3F4_F5D5PHI1X1_wr_en),
.number_out(CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5_number),
.read_add(CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5_read_add),
.data_out(CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5),
.start(ME_F3F4_F5D5PHI1X1_start),
.done(CM_F3F4_F5D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F5D5PHI1X2_CM_F3F4_F5D5PHI1X2;
wire ME_F3F4_F5D5PHI1X2_CM_F3F4_F5D5PHI1X2_wr_en;
wire [5:0] CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5_number;
wire [8:0] CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5_read_add;
wire [11:0] CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5;
CandidateMatch  CM_F3F4_F5D5PHI1X2(
.data_in(ME_F3F4_F5D5PHI1X2_CM_F3F4_F5D5PHI1X2),
.enable(ME_F3F4_F5D5PHI1X2_CM_F3F4_F5D5PHI1X2_wr_en),
.number_out(CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5_number),
.read_add(CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5_read_add),
.data_out(CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5),
.start(ME_F3F4_F5D5PHI1X2_start),
.done(CM_F3F4_F5D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F5D5PHI2X1_CM_F3F4_F5D5PHI2X1;
wire ME_F3F4_F5D5PHI2X1_CM_F3F4_F5D5PHI2X1_wr_en;
wire [5:0] CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5_number;
wire [8:0] CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5_read_add;
wire [11:0] CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5;
CandidateMatch  CM_F3F4_F5D5PHI2X1(
.data_in(ME_F3F4_F5D5PHI2X1_CM_F3F4_F5D5PHI2X1),
.enable(ME_F3F4_F5D5PHI2X1_CM_F3F4_F5D5PHI2X1_wr_en),
.number_out(CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5_number),
.read_add(CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5_read_add),
.data_out(CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5),
.start(ME_F3F4_F5D5PHI2X1_start),
.done(CM_F3F4_F5D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F5D5PHI2X2_CM_F3F4_F5D5PHI2X2;
wire ME_F3F4_F5D5PHI2X2_CM_F3F4_F5D5PHI2X2_wr_en;
wire [5:0] CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5_number;
wire [8:0] CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5_read_add;
wire [11:0] CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5;
CandidateMatch  CM_F3F4_F5D5PHI2X2(
.data_in(ME_F3F4_F5D5PHI2X2_CM_F3F4_F5D5PHI2X2),
.enable(ME_F3F4_F5D5PHI2X2_CM_F3F4_F5D5PHI2X2_wr_en),
.number_out(CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5_number),
.read_add(CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5_read_add),
.data_out(CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5),
.start(ME_F3F4_F5D5PHI2X2_start),
.done(CM_F3F4_F5D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F5D5PHI3X1_CM_F3F4_F5D5PHI3X1;
wire ME_F3F4_F5D5PHI3X1_CM_F3F4_F5D5PHI3X1_wr_en;
wire [5:0] CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5_number;
wire [8:0] CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5_read_add;
wire [11:0] CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5;
CandidateMatch  CM_F3F4_F5D5PHI3X1(
.data_in(ME_F3F4_F5D5PHI3X1_CM_F3F4_F5D5PHI3X1),
.enable(ME_F3F4_F5D5PHI3X1_CM_F3F4_F5D5PHI3X1_wr_en),
.number_out(CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5_number),
.read_add(CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5_read_add),
.data_out(CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5),
.start(ME_F3F4_F5D5PHI3X1_start),
.done(CM_F3F4_F5D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F5D5PHI3X2_CM_F3F4_F5D5PHI3X2;
wire ME_F3F4_F5D5PHI3X2_CM_F3F4_F5D5PHI3X2_wr_en;
wire [5:0] CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5_number;
wire [8:0] CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5_read_add;
wire [11:0] CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5;
CandidateMatch  CM_F3F4_F5D5PHI3X2(
.data_in(ME_F3F4_F5D5PHI3X2_CM_F3F4_F5D5PHI3X2),
.enable(ME_F3F4_F5D5PHI3X2_CM_F3F4_F5D5PHI3X2_wr_en),
.number_out(CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5_number),
.read_add(CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5_read_add),
.data_out(CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5),
.start(ME_F3F4_F5D5PHI3X2_start),
.done(CM_F3F4_F5D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F5D5PHI4X1_CM_F3F4_F5D5PHI4X1;
wire ME_F3F4_F5D5PHI4X1_CM_F3F4_F5D5PHI4X1_wr_en;
wire [5:0] CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5_number;
wire [8:0] CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5_read_add;
wire [11:0] CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5;
CandidateMatch  CM_F3F4_F5D5PHI4X1(
.data_in(ME_F3F4_F5D5PHI4X1_CM_F3F4_F5D5PHI4X1),
.enable(ME_F3F4_F5D5PHI4X1_CM_F3F4_F5D5PHI4X1_wr_en),
.number_out(CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5_number),
.read_add(CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5_read_add),
.data_out(CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5),
.start(ME_F3F4_F5D5PHI4X1_start),
.done(CM_F3F4_F5D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_F3F4_F5D5PHI4X2_CM_F3F4_F5D5PHI4X2;
wire ME_F3F4_F5D5PHI4X2_CM_F3F4_F5D5PHI4X2_wr_en;
wire [5:0] CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5_number;
wire [8:0] CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5_read_add;
wire [11:0] CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5;
CandidateMatch  CM_F3F4_F5D5PHI4X2(
.data_in(ME_F3F4_F5D5PHI4X2_CM_F3F4_F5D5PHI4X2),
.enable(ME_F3F4_F5D5PHI4X2_CM_F3F4_F5D5PHI4X2_wr_en),
.number_out(CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5_number),
.read_add(CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5_read_add),
.data_out(CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5),
.start(ME_F3F4_F5D5PHI4X2_start),
.done(CM_F3F4_F5D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PRD_F5D5_F3F4_AP_F3F4_F5D5;
wire PRD_F5D5_F3F4_AP_F3F4_F5D5_wr_en;
wire [8:0] AP_F3F4_F5D5_MC_F3F4_F5D5_read_add;
wire [55:0] AP_F3F4_F5D5_MC_F3F4_F5D5;
AllProj #(1'b0,1'b1) AP_F3F4_F5D5(
.data_in(PRD_F5D5_F3F4_AP_F3F4_F5D5),
.enable(PRD_F5D5_F3F4_AP_F3F4_F5D5_wr_en),
.read_add(AP_F3F4_F5D5_MC_F3F4_F5D5_read_add),
.data_out(AP_F3F4_F5D5_MC_F3F4_F5D5),
.start(PRD_F5D5_F3F4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMRD_F5D5_AS_F5D5n2;
wire VMRD_F5D5_AS_F5D5n2_wr_en;
wire [10:0] AS_F5D5n2_MC_F3F4_F5D5_read_add;
wire [35:0] AS_F5D5n2_MC_F3F4_F5D5;
AllStubs  AS_F5D5n2(
.data_in(VMRD_F5D5_AS_F5D5n2),
.enable(VMRD_F5D5_AS_F5D5n2_wr_en),
.read_add_MC(AS_F5D5n2_MC_F3F4_F5D5_read_add),
.data_out_MC(AS_F5D5n2_MC_F3F4_F5D5),
.start(VMRD_F5D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F3D5_FM_F1F2_F3D5_ToMinus;
wire MC_F1F2_F3D5_FM_F1F2_F3D5_ToMinus_wr_en;
wire [5:0] FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus_number;
wire [9:0] FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus_read_add;
wire [39:0] FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus;
FullMatch #(128) FM_F1F2_F3D5_ToMinus(
.data_in(MC_F1F2_F3D5_FM_F1F2_F3D5_ToMinus),
.enable(MC_F1F2_F3D5_FM_F1F2_F3D5_ToMinus_wr_en),
.number_out(FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus_number),
.read_add(FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus_read_add),
.data_out(FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus),
.read_en(1'b1),
.start(MC_F1F2_F3D5_start),
.done(FM_F1F2_F3D5_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F4D5_FM_F1F2_F4D5_ToMinus;
wire MC_F1F2_F4D5_FM_F1F2_F4D5_ToMinus_wr_en;
wire [5:0] FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus_number;
wire [9:0] FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus_read_add;
wire [39:0] FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus;
FullMatch #(128) FM_F1F2_F4D5_ToMinus(
.data_in(MC_F1F2_F4D5_FM_F1F2_F4D5_ToMinus),
.enable(MC_F1F2_F4D5_FM_F1F2_F4D5_ToMinus_wr_en),
.number_out(FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus_number),
.read_add(FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus_read_add),
.data_out(FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus),
.read_en(1'b1),
.start(MC_F1F2_F4D5_start),
.done(FM_F1F2_F4D5_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F5D5_FM_F1F2_F5D5_ToMinus;
wire MC_F1F2_F5D5_FM_F1F2_F5D5_ToMinus_wr_en;
wire [5:0] FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus_number;
wire [9:0] FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus_read_add;
wire [39:0] FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus;
FullMatch #(128) FM_F1F2_F5D5_ToMinus(
.data_in(MC_F1F2_F5D5_FM_F1F2_F5D5_ToMinus),
.enable(MC_F1F2_F5D5_FM_F1F2_F5D5_ToMinus_wr_en),
.number_out(FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus_number),
.read_add(FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus_read_add),
.data_out(FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus),
.read_en(1'b1),
.start(MC_F1F2_F5D5_start),
.done(FM_F1F2_F5D5_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToMinus;
wire MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToMinus_wr_en;
wire [5:0] FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus_number;
wire [9:0] FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus_read_add;
wire [39:0] FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus;
FullMatch #(128) FM_FL3FL4_F1D5_ToMinus(
.data_in(MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToMinus),
.enable(MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToMinus_wr_en),
.number_out(FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus_number),
.read_add(FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus_read_add),
.data_out(FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus),
.read_en(1'b1),
.start(MC_F3F4_F1D5_start),
.done(FM_FL3FL4_F1D5_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToMinus;
wire MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToMinus_wr_en;
wire [5:0] FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus_number;
wire [9:0] FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus_read_add;
wire [39:0] FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus;
FullMatch #(128) FM_FL3FL4_F2D5_ToMinus(
.data_in(MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToMinus),
.enable(MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToMinus_wr_en),
.number_out(FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus_number),
.read_add(FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus_read_add),
.data_out(FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus),
.read_en(1'b1),
.start(MC_F3F4_F2D5_start),
.done(FM_FL3FL4_F2D5_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F5D5_FM_F3F4_F5D5_ToMinus;
wire MC_F3F4_F5D5_FM_F3F4_F5D5_ToMinus_wr_en;
wire [5:0] FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus_number;
wire [9:0] FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus_read_add;
wire [39:0] FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus;
FullMatch #(128) FM_F3F4_F5D5_ToMinus(
.data_in(MC_F3F4_F5D5_FM_F3F4_F5D5_ToMinus),
.enable(MC_F3F4_F5D5_FM_F3F4_F5D5_ToMinus_wr_en),
.number_out(FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus_number),
.read_add(FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus_read_add),
.data_out(FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus),
.read_en(1'b1),
.start(MC_F3F4_F5D5_start),
.done(FM_F3F4_F5D5_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F3D5_FM_F1F2_F3D5_ToPlus;
wire MC_F1F2_F3D5_FM_F1F2_F3D5_ToPlus_wr_en;
wire [5:0] FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus_number;
wire [9:0] FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus_read_add;
wire [39:0] FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus;
FullMatch #(128) FM_F1F2_F3D5_ToPlus(
.data_in(MC_F1F2_F3D5_FM_F1F2_F3D5_ToPlus),
.enable(MC_F1F2_F3D5_FM_F1F2_F3D5_ToPlus_wr_en),
.number_out(FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus_number),
.read_add(FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus_read_add),
.data_out(FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus),
.read_en(1'b1),
.start(MC_F1F2_F3D5_start),
.done(FM_F1F2_F3D5_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F4D5_FM_F1F2_F4D5_ToPlus;
wire MC_F1F2_F4D5_FM_F1F2_F4D5_ToPlus_wr_en;
wire [5:0] FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus_number;
wire [9:0] FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus_read_add;
wire [39:0] FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus;
FullMatch #(128) FM_F1F2_F4D5_ToPlus(
.data_in(MC_F1F2_F4D5_FM_F1F2_F4D5_ToPlus),
.enable(MC_F1F2_F4D5_FM_F1F2_F4D5_ToPlus_wr_en),
.number_out(FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus_number),
.read_add(FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus_read_add),
.data_out(FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus),
.read_en(1'b1),
.start(MC_F1F2_F4D5_start),
.done(FM_F1F2_F4D5_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F5D5_FM_F1F2_F5D5_ToPlus;
wire MC_F1F2_F5D5_FM_F1F2_F5D5_ToPlus_wr_en;
wire [5:0] FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus_number;
wire [9:0] FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus_read_add;
wire [39:0] FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus;
FullMatch #(128) FM_F1F2_F5D5_ToPlus(
.data_in(MC_F1F2_F5D5_FM_F1F2_F5D5_ToPlus),
.enable(MC_F1F2_F5D5_FM_F1F2_F5D5_ToPlus_wr_en),
.number_out(FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus_number),
.read_add(FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus_read_add),
.data_out(FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus),
.read_en(1'b1),
.start(MC_F1F2_F5D5_start),
.done(FM_F1F2_F5D5_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToPlus;
wire MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToPlus_wr_en;
wire [5:0] FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus_number;
wire [9:0] FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus_read_add;
wire [39:0] FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus;
FullMatch #(128) FM_FL3FL4_F1D5_ToPlus(
.data_in(MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToPlus),
.enable(MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToPlus_wr_en),
.number_out(FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus_number),
.read_add(FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus_read_add),
.data_out(FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus),
.read_en(1'b1),
.start(MC_F3F4_F1D5_start),
.done(FM_FL3FL4_F1D5_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToPlus;
wire MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToPlus_wr_en;
wire [5:0] FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus_number;
wire [9:0] FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus_read_add;
wire [39:0] FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus;
FullMatch #(128) FM_FL3FL4_F2D5_ToPlus(
.data_in(MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToPlus),
.enable(MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToPlus_wr_en),
.number_out(FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus_number),
.read_add(FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus_read_add),
.data_out(FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus),
.read_en(1'b1),
.start(MC_F3F4_F2D5_start),
.done(FM_FL3FL4_F2D5_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F5D5_FM_F3F4_F5D5_ToPlus;
wire MC_F3F4_F5D5_FM_F3F4_F5D5_ToPlus_wr_en;
wire [5:0] FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus_number;
wire [9:0] FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus_read_add;
wire [39:0] FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus;
FullMatch #(128) FM_F3F4_F5D5_ToPlus(
.data_in(MC_F3F4_F5D5_FM_F3F4_F5D5_ToPlus),
.enable(MC_F3F4_F5D5_FM_F3F4_F5D5_ToPlus_wr_en),
.number_out(FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus_number),
.read_add(FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus_read_add),
.data_out(FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus),
.read_en(1'b1),
.start(MC_F3F4_F5D5_start),
.done(FM_F3F4_F5D5_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F3D5_FM_F1F2_F3D5;
wire MC_F1F2_F3D5_FM_F1F2_F3D5_wr_en;
wire [5:0] FM_F1F2_F3D5_FT_F1F2_number;
wire [9:0] FM_F1F2_F3D5_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F3D5_FT_F1F2;
wire FM_F1F2_F3D5_FT_F1F2_read_en;
FullMatch  FM_F1F2_F3D5(
.data_in(MC_F1F2_F3D5_FM_F1F2_F3D5),
.enable(MC_F1F2_F3D5_FM_F1F2_F3D5_wr_en),
.number_out(FM_F1F2_F3D5_FT_F1F2_number),
.read_add(FM_F1F2_F3D5_FT_F1F2_read_add),
.data_out(FM_F1F2_F3D5_FT_F1F2),
.read_en(FM_F1F2_F3D5_FT_F1F2_read_en),
.start(MC_F1F2_F3D5_start),
.done(FM_F1F2_F3D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F4D5_FM_F1F2_F4D5;
wire MC_F1F2_F4D5_FM_F1F2_F4D5_wr_en;
wire [5:0] FM_F1F2_F4D5_FT_F1F2_number;
wire [9:0] FM_F1F2_F4D5_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F4D5_FT_F1F2;
wire FM_F1F2_F4D5_FT_F1F2_read_en;
FullMatch  FM_F1F2_F4D5(
.data_in(MC_F1F2_F4D5_FM_F1F2_F4D5),
.enable(MC_F1F2_F4D5_FM_F1F2_F4D5_wr_en),
.number_out(FM_F1F2_F4D5_FT_F1F2_number),
.read_add(FM_F1F2_F4D5_FT_F1F2_read_add),
.data_out(FM_F1F2_F4D5_FT_F1F2),
.read_en(FM_F1F2_F4D5_FT_F1F2_read_en),
.start(MC_F1F2_F4D5_start),
.done(FM_F1F2_F4D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F1F2_F5D5_FM_F1F2_F5D5;
wire MC_F1F2_F5D5_FM_F1F2_F5D5_wr_en;
wire [5:0] FM_F1F2_F5D5_FT_F1F2_number;
wire [9:0] FM_F1F2_F5D5_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F5D5_FT_F1F2;
wire FM_F1F2_F5D5_FT_F1F2_read_en;
FullMatch  FM_F1F2_F5D5(
.data_in(MC_F1F2_F5D5_FM_F1F2_F5D5),
.enable(MC_F1F2_F5D5_FM_F1F2_F5D5_wr_en),
.number_out(FM_F1F2_F5D5_FT_F1F2_number),
.read_add(FM_F1F2_F5D5_FT_F1F2_read_add),
.data_out(FM_F1F2_F5D5_FT_F1F2),
.read_en(FM_F1F2_F5D5_FT_F1F2_read_en),
.start(MC_F1F2_F5D5_start),
.done(FM_F1F2_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_F1D5F2D5_TPAR_F1D5F2D5;
wire TC_F1D5F2D5_TPAR_F1D5F2D5_wr_en;
wire [10:0] TPAR_F1D5F2D5_FT_F1F2_read_add;
wire [67:0] TPAR_F1D5F2D5_FT_F1F2;
TrackletParameters  TPAR_F1D5F2D5(
.data_in(TC_F1D5F2D5_TPAR_F1D5F2D5),
.enable(TC_F1D5F2D5_TPAR_F1D5F2D5_wr_en),
.read_add(TPAR_F1D5F2D5_FT_F1F2_read_add),
.data_out(TPAR_F1D5F2D5_FT_F1F2),
.start(TC_F1D5F2D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Minus_FM_F1F2_F3_FromMinus;
wire MT_FDSK_Minus_FM_F1F2_F3_FromMinus_wr_en;
wire [5:0] FM_F1F2_F3_FromMinus_FT_F1F2_number;
wire [9:0] FM_F1F2_F3_FromMinus_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F3_FromMinus_FT_F1F2;
wire FM_F1F2_F3_FromMinus_FT_F1F2_read_en;
FullMatch #(128) FM_F1F2_F3_FromMinus(
.data_in(MT_FDSK_Minus_FM_F1F2_F3_FromMinus),
.enable(MT_FDSK_Minus_FM_F1F2_F3_FromMinus_wr_en),
.number_out(FM_F1F2_F3_FromMinus_FT_F1F2_number),
.read_add(FM_F1F2_F3_FromMinus_FT_F1F2_read_add),
.data_out(FM_F1F2_F3_FromMinus_FT_F1F2),
.read_en(FM_F1F2_F3_FromMinus_FT_F1F2_read_en),
.start(MT_FDSK_Minus_start),
.done(FM_F1F2_F3_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Minus_FM_F1F2_F4_FromMinus;
wire MT_FDSK_Minus_FM_F1F2_F4_FromMinus_wr_en;
wire [5:0] FM_F1F2_F4_FromMinus_FT_F1F2_number;
wire [9:0] FM_F1F2_F4_FromMinus_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F4_FromMinus_FT_F1F2;
wire FM_F1F2_F4_FromMinus_FT_F1F2_read_en;
FullMatch #(128) FM_F1F2_F4_FromMinus(
.data_in(MT_FDSK_Minus_FM_F1F2_F4_FromMinus),
.enable(MT_FDSK_Minus_FM_F1F2_F4_FromMinus_wr_en),
.number_out(FM_F1F2_F4_FromMinus_FT_F1F2_number),
.read_add(FM_F1F2_F4_FromMinus_FT_F1F2_read_add),
.data_out(FM_F1F2_F4_FromMinus_FT_F1F2),
.read_en(FM_F1F2_F4_FromMinus_FT_F1F2_read_en),
.start(MT_FDSK_Minus_start),
.done(FM_F1F2_F4_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Minus_FM_F1F2_F5_FromMinus;
wire MT_FDSK_Minus_FM_F1F2_F5_FromMinus_wr_en;
wire [5:0] FM_F1F2_F5_FromMinus_FT_F1F2_number;
wire [9:0] FM_F1F2_F5_FromMinus_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F5_FromMinus_FT_F1F2;
wire FM_F1F2_F5_FromMinus_FT_F1F2_read_en;
FullMatch #(128) FM_F1F2_F5_FromMinus(
.data_in(MT_FDSK_Minus_FM_F1F2_F5_FromMinus),
.enable(MT_FDSK_Minus_FM_F1F2_F5_FromMinus_wr_en),
.number_out(FM_F1F2_F5_FromMinus_FT_F1F2_number),
.read_add(FM_F1F2_F5_FromMinus_FT_F1F2_read_add),
.data_out(FM_F1F2_F5_FromMinus_FT_F1F2),
.read_en(FM_F1F2_F5_FromMinus_FT_F1F2_read_en),
.start(MT_FDSK_Minus_start),
.done(FM_F1F2_F5_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Plus_FM_F1F2_F3_FromPlus;
wire MT_FDSK_Plus_FM_F1F2_F3_FromPlus_wr_en;
wire [5:0] FM_F1F2_F3_FromPlus_FT_F1F2_number;
wire [9:0] FM_F1F2_F3_FromPlus_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F3_FromPlus_FT_F1F2;
wire FM_F1F2_F3_FromPlus_FT_F1F2_read_en;
FullMatch #(128) FM_F1F2_F3_FromPlus(
.data_in(MT_FDSK_Plus_FM_F1F2_F3_FromPlus),
.enable(MT_FDSK_Plus_FM_F1F2_F3_FromPlus_wr_en),
.number_out(FM_F1F2_F3_FromPlus_FT_F1F2_number),
.read_add(FM_F1F2_F3_FromPlus_FT_F1F2_read_add),
.data_out(FM_F1F2_F3_FromPlus_FT_F1F2),
.read_en(FM_F1F2_F3_FromPlus_FT_F1F2_read_en),
.start(MT_FDSK_Plus_start),
.done(FM_F1F2_F3_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Plus_FM_F1F2_F4_FromPlus;
wire MT_FDSK_Plus_FM_F1F2_F4_FromPlus_wr_en;
wire [5:0] FM_F1F2_F4_FromPlus_FT_F1F2_number;
wire [9:0] FM_F1F2_F4_FromPlus_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F4_FromPlus_FT_F1F2;
wire FM_F1F2_F4_FromPlus_FT_F1F2_read_en;
FullMatch #(128) FM_F1F2_F4_FromPlus(
.data_in(MT_FDSK_Plus_FM_F1F2_F4_FromPlus),
.enable(MT_FDSK_Plus_FM_F1F2_F4_FromPlus_wr_en),
.number_out(FM_F1F2_F4_FromPlus_FT_F1F2_number),
.read_add(FM_F1F2_F4_FromPlus_FT_F1F2_read_add),
.data_out(FM_F1F2_F4_FromPlus_FT_F1F2),
.read_en(FM_F1F2_F4_FromPlus_FT_F1F2_read_en),
.start(MT_FDSK_Plus_start),
.done(FM_F1F2_F4_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Plus_FM_F1F2_F5_FromPlus;
wire MT_FDSK_Plus_FM_F1F2_F5_FromPlus_wr_en;
wire [5:0] FM_F1F2_F5_FromPlus_FT_F1F2_number;
wire [9:0] FM_F1F2_F5_FromPlus_FT_F1F2_read_add;
wire [39:0] FM_F1F2_F5_FromPlus_FT_F1F2;
wire FM_F1F2_F5_FromPlus_FT_F1F2_read_en;
FullMatch #(128) FM_F1F2_F5_FromPlus(
.data_in(MT_FDSK_Plus_FM_F1F2_F5_FromPlus),
.enable(MT_FDSK_Plus_FM_F1F2_F5_FromPlus_wr_en),
.number_out(FM_F1F2_F5_FromPlus_FT_F1F2_number),
.read_add(FM_F1F2_F5_FromPlus_FT_F1F2_read_add),
.data_out(FM_F1F2_F5_FromPlus_FT_F1F2),
.read_en(FM_F1F2_F5_FromPlus_FT_F1F2_read_en),
.start(MT_FDSK_Plus_start),
.done(FM_F1F2_F5_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F1D5_FM_F3F4_F1D5;
wire MC_F3F4_F1D5_FM_F3F4_F1D5_wr_en;
wire [5:0] FM_F3F4_F1D5_FT_F3F4_number;
wire [9:0] FM_F3F4_F1D5_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F1D5_FT_F3F4;
wire FM_F3F4_F1D5_FT_F3F4_read_en;
FullMatch  FM_F3F4_F1D5(
.data_in(MC_F3F4_F1D5_FM_F3F4_F1D5),
.enable(MC_F3F4_F1D5_FM_F3F4_F1D5_wr_en),
.number_out(FM_F3F4_F1D5_FT_F3F4_number),
.read_add(FM_F3F4_F1D5_FT_F3F4_read_add),
.data_out(FM_F3F4_F1D5_FT_F3F4),
.read_en(FM_F3F4_F1D5_FT_F3F4_read_en),
.start(MC_F3F4_F1D5_start),
.done(FM_F3F4_F1D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F2D5_FM_F3F4_F2D5;
wire MC_F3F4_F2D5_FM_F3F4_F2D5_wr_en;
wire [5:0] FM_F3F4_F2D5_FT_F3F4_number;
wire [9:0] FM_F3F4_F2D5_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F2D5_FT_F3F4;
wire FM_F3F4_F2D5_FT_F3F4_read_en;
FullMatch  FM_F3F4_F2D5(
.data_in(MC_F3F4_F2D5_FM_F3F4_F2D5),
.enable(MC_F3F4_F2D5_FM_F3F4_F2D5_wr_en),
.number_out(FM_F3F4_F2D5_FT_F3F4_number),
.read_add(FM_F3F4_F2D5_FT_F3F4_read_add),
.data_out(FM_F3F4_F2D5_FT_F3F4),
.read_en(FM_F3F4_F2D5_FT_F3F4_read_en),
.start(MC_F3F4_F2D5_start),
.done(FM_F3F4_F2D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_F3F4_F5D5_FM_F3F4_F5D5;
wire MC_F3F4_F5D5_FM_F3F4_F5D5_wr_en;
wire [5:0] FM_F3F4_F5D5_FT_F3F4_number;
wire [9:0] FM_F3F4_F5D5_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F5D5_FT_F3F4;
wire FM_F3F4_F5D5_FT_F3F4_read_en;
FullMatch  FM_F3F4_F5D5(
.data_in(MC_F3F4_F5D5_FM_F3F4_F5D5),
.enable(MC_F3F4_F5D5_FM_F3F4_F5D5_wr_en),
.number_out(FM_F3F4_F5D5_FT_F3F4_number),
.read_add(FM_F3F4_F5D5_FT_F3F4_read_add),
.data_out(FM_F3F4_F5D5_FT_F3F4),
.read_en(FM_F3F4_F5D5_FT_F3F4_read_en),
.start(MC_F3F4_F5D5_start),
.done(FM_F3F4_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_F3D5F4D5_TPAR_F3D5F4D5;
wire TC_F3D5F4D5_TPAR_F3D5F4D5_wr_en;
wire [10:0] TPAR_F3D5F4D5_FT_F3F4_read_add;
wire [67:0] TPAR_F3D5F4D5_FT_F3F4;
TrackletParameters  TPAR_F3D5F4D5(
.data_in(TC_F3D5F4D5_TPAR_F3D5F4D5),
.enable(TC_F3D5F4D5_TPAR_F3D5F4D5_wr_en),
.read_add(TPAR_F3D5F4D5_FT_F3F4_read_add),
.data_out(TPAR_F3D5F4D5_FT_F3F4),
.start(TC_F3D5F4D5_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Minus_FM_F3F4_F1_FromMinus;
wire MT_FDSK_Minus_FM_F3F4_F1_FromMinus_wr_en;
wire [5:0] FM_F3F4_F1_FromMinus_FT_F3F4_number;
wire [9:0] FM_F3F4_F1_FromMinus_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F1_FromMinus_FT_F3F4;
wire FM_F3F4_F1_FromMinus_FT_F3F4_read_en;
FullMatch #(128) FM_F3F4_F1_FromMinus(
.data_in(MT_FDSK_Minus_FM_F3F4_F1_FromMinus),
.enable(MT_FDSK_Minus_FM_F3F4_F1_FromMinus_wr_en),
.number_out(FM_F3F4_F1_FromMinus_FT_F3F4_number),
.read_add(FM_F3F4_F1_FromMinus_FT_F3F4_read_add),
.data_out(FM_F3F4_F1_FromMinus_FT_F3F4),
.read_en(FM_F3F4_F1_FromMinus_FT_F3F4_read_en),
.start(MT_FDSK_Minus_start),
.done(FM_F3F4_F1_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Minus_FM_F3F4_F2_FromMinus;
wire MT_FDSK_Minus_FM_F3F4_F2_FromMinus_wr_en;
wire [5:0] FM_F3F4_F2_FromMinus_FT_F3F4_number;
wire [9:0] FM_F3F4_F2_FromMinus_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F2_FromMinus_FT_F3F4;
wire FM_F3F4_F2_FromMinus_FT_F3F4_read_en;
FullMatch #(128) FM_F3F4_F2_FromMinus(
.data_in(MT_FDSK_Minus_FM_F3F4_F2_FromMinus),
.enable(MT_FDSK_Minus_FM_F3F4_F2_FromMinus_wr_en),
.number_out(FM_F3F4_F2_FromMinus_FT_F3F4_number),
.read_add(FM_F3F4_F2_FromMinus_FT_F3F4_read_add),
.data_out(FM_F3F4_F2_FromMinus_FT_F3F4),
.read_en(FM_F3F4_F2_FromMinus_FT_F3F4_read_en),
.start(MT_FDSK_Minus_start),
.done(FM_F3F4_F2_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Minus_FM_F3F4_F5_FromMinus;
wire MT_FDSK_Minus_FM_F3F4_F5_FromMinus_wr_en;
wire [5:0] FM_F3F4_F5_FromMinus_FT_F3F4_number;
wire [9:0] FM_F3F4_F5_FromMinus_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F5_FromMinus_FT_F3F4;
wire FM_F3F4_F5_FromMinus_FT_F3F4_read_en;
FullMatch #(128) FM_F3F4_F5_FromMinus(
.data_in(MT_FDSK_Minus_FM_F3F4_F5_FromMinus),
.enable(MT_FDSK_Minus_FM_F3F4_F5_FromMinus_wr_en),
.number_out(FM_F3F4_F5_FromMinus_FT_F3F4_number),
.read_add(FM_F3F4_F5_FromMinus_FT_F3F4_read_add),
.data_out(FM_F3F4_F5_FromMinus_FT_F3F4),
.read_en(FM_F3F4_F5_FromMinus_FT_F3F4_read_en),
.start(MT_FDSK_Minus_start),
.done(FM_F3F4_F5_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Plus_FM_F3F4_F1_FromPlus;
wire MT_FDSK_Plus_FM_F3F4_F1_FromPlus_wr_en;
wire [5:0] FM_F3F4_F1_FromPlus_FT_F3F4_number;
wire [9:0] FM_F3F4_F1_FromPlus_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F1_FromPlus_FT_F3F4;
wire FM_F3F4_F1_FromPlus_FT_F3F4_read_en;
FullMatch #(128) FM_F3F4_F1_FromPlus(
.data_in(MT_FDSK_Plus_FM_F3F4_F1_FromPlus),
.enable(MT_FDSK_Plus_FM_F3F4_F1_FromPlus_wr_en),
.number_out(FM_F3F4_F1_FromPlus_FT_F3F4_number),
.read_add(FM_F3F4_F1_FromPlus_FT_F3F4_read_add),
.data_out(FM_F3F4_F1_FromPlus_FT_F3F4),
.read_en(FM_F3F4_F1_FromPlus_FT_F3F4_read_en),
.start(MT_FDSK_Plus_start),
.done(FM_F3F4_F1_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Plus_FM_F3F4_F2_FromPlus;
wire MT_FDSK_Plus_FM_F3F4_F2_FromPlus_wr_en;
wire [5:0] FM_F3F4_F2_FromPlus_FT_F3F4_number;
wire [9:0] FM_F3F4_F2_FromPlus_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F2_FromPlus_FT_F3F4;
wire FM_F3F4_F2_FromPlus_FT_F3F4_read_en;
FullMatch #(128) FM_F3F4_F2_FromPlus(
.data_in(MT_FDSK_Plus_FM_F3F4_F2_FromPlus),
.enable(MT_FDSK_Plus_FM_F3F4_F2_FromPlus_wr_en),
.number_out(FM_F3F4_F2_FromPlus_FT_F3F4_number),
.read_add(FM_F3F4_F2_FromPlus_FT_F3F4_read_add),
.data_out(FM_F3F4_F2_FromPlus_FT_F3F4),
.read_en(FM_F3F4_F2_FromPlus_FT_F3F4_read_en),
.start(MT_FDSK_Plus_start),
.done(FM_F3F4_F2_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_FDSK_Plus_FM_F3F4_F5_FromPlus;
wire MT_FDSK_Plus_FM_F3F4_F5_FromPlus_wr_en;
wire [5:0] FM_F3F4_F5_FromPlus_FT_F3F4_number;
wire [9:0] FM_F3F4_F5_FromPlus_FT_F3F4_read_add;
wire [39:0] FM_F3F4_F5_FromPlus_FT_F3F4;
wire FM_F3F4_F5_FromPlus_FT_F3F4_read_en;
FullMatch #(128) FM_F3F4_F5_FromPlus(
.data_in(MT_FDSK_Plus_FM_F3F4_F5_FromPlus),
.enable(MT_FDSK_Plus_FM_F3F4_F5_FromPlus_wr_en),
.number_out(FM_F3F4_F5_FromPlus_FT_F3F4_number),
.read_add(FM_F3F4_F5_FromPlus_FT_F3F4_read_add),
.data_out(FM_F3F4_F5_FromPlus_FT_F3F4),
.read_en(FM_F3F4_F5_FromPlus_FT_F3F4_read_en),
.start(MT_FDSK_Plus_start),
.done(FM_F3F4_F5_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] FT_F1F2_TF_F1F2;
wire FT_F1F2_TF_F1F2_wr_en;
wire [8:0] TF_F1F2_PD_read_add;
wire [125:0] TF_F1F2_PD;
TrackFit  TF_F1F2(
.data_in(FT_F1F2_TF_F1F2),
.enable(FT_F1F2_TF_F1F2_wr_en),
.read_add(TF_F1F2_PD_read_add),
.data_out(TF_F1F2_PD),
.start(FT_F1F2_start),
.done(TF_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] FT_F3F4_TF_F3F4;
wire FT_F3F4_TF_F3F4_wr_en;
wire [8:0] TF_F3F4_PD_read_add;
wire [125:0] TF_F3F4_PD;
TrackFit  TF_F3F4(
.data_in(FT_F3F4_TF_F3F4),
.enable(FT_F3F4_TF_F3F4_wr_en),
.read_add(TF_F3F4_PD_read_add),
.data_out(TF_F3F4_PD),
.start(FT_F3F4_start),
.done(TF_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] PD_CT_F1F2;
wire PD_CT_F1F2_wr_en;
//wire CT_F1F2_DataStream;
CleanTrack  CT_F1F2(
.data_in(PD_CT_F1F2),
.enable(PD_CT_F1F2_wr_en),
.data_out(CT_F1F2_DataStream),
.start(PD_start),
.done(CT_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] PD_CT_F3F4;
wire PD_CT_F3F4_wr_en;
//wire CT_F3F4_DataStream;
CleanTrack  CT_F3F4(
.data_in(PD_CT_F3F4),
.enable(PD_CT_F3F4_wr_en),
.data_out(CT_F3F4_DataStream),
.start(PD_start),
.done(CT_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L3F3F5") PT_L3F3F5_Plus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus_number),
.read_add_projin_disk_2(TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus_read_add),
.projin_disk_2(TPROJ_ToPlus_F1D5F2D5_F5_PT_L3F3F5_Plus),
.number_in_projin_disk_3(TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus_number),
.read_add_projin_disk_3(TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus_read_add),
.projin_disk_3(TPROJ_ToPlus_F3D5F4D5_F5_PT_L3F3F5_Plus),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus_number),
.read_add_projin_disk_7(TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus_read_add),
.projin_disk_7(TPROJ_ToPlus_F1D5F2D5_F3_PT_L3F3F5_Plus),
.number_in_projin_disk_8(6'b0),
.number_in_projin_disk_9(6'b0),
.number_in_projin_layer_1(6'b0),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(6'b0),
.number_in_projin_layer_5(6'b0),
.number_in_projin_layer_6(6'b0),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L3F3F5_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L3F3F5_Plus_From_DataStream),
.projout_disk_1(PT_L3F3F5_Plus_TPROJ_FromPlus_F3D5_F1F2),
.valid_disk_1(PT_L3F3F5_Plus_TPROJ_FromPlus_F3D5_F1F2_wr_en),
.projout_disk_3(PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F1F2),
.valid_disk_3(PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F1F2_wr_en),
.projout_disk_5(PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F3F4),
.valid_disk_5(PT_L3F3F5_Plus_TPROJ_FromPlus_F5D5_F3F4_wr_en),
.valid_proj_data_stream(PT_L3F3F5_Plus_To_DataStream_en),
.proj_data_stream(PT_L3F3F5_Plus_To_DataStream),
.start(TPROJ_ToPlus_F1D5F2D5_F5_start),
.done(PT_L3F3F5_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L2L4F2") PT_L2L4F2_Plus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus_number),
.read_add_projin_disk_2(TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus_read_add),
.projin_disk_2(TPROJ_ToPlus_F3D5F4D5_F2_PT_L2L4F2_Plus),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_disk_8(6'b0),
.number_in_projin_disk_9(6'b0),
.number_in_projin_layer_1(6'b0),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(6'b0),
.number_in_projin_layer_5(6'b0),
.number_in_projin_layer_6(6'b0),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L2L4F2_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L2L4F2_Plus_From_DataStream),
.projout_disk_1(PT_L2L4F2_Plus_TPROJ_FromPlus_F2D5_F3F4),
.valid_disk_1(PT_L2L4F2_Plus_TPROJ_FromPlus_F2D5_F3F4_wr_en),
.valid_proj_data_stream(PT_L2L4F2_Plus_To_DataStream_en),
.proj_data_stream(PT_L2L4F2_Plus_To_DataStream),
.start(TPROJ_ToPlus_F3D5F4D5_F2_start),
.done(PT_L2L4F2_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("F1L5") PT_F1L5_Plus(
.number_in_projin_disk_1(TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus_number),
.read_add_projin_disk_1(TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus_read_add),
.projin_disk_1(TPROJ_ToPlus_F3D5F4D5_F1_PT_F1L5_Plus),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_disk_8(6'b0),
.number_in_projin_disk_9(6'b0),
.number_in_projin_layer_1(6'b0),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(6'b0),
.number_in_projin_layer_5(6'b0),
.number_in_projin_layer_6(6'b0),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_F1L5_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_F1L5_Plus_From_DataStream),
.projout_disk_1(PT_F1L5_Plus_TPROJ_FromPlus_F1D5_F3F4),
.valid_disk_1(PT_F1L5_Plus_TPROJ_FromPlus_F1D5_F3F4_wr_en),
.valid_proj_data_stream(PT_F1L5_Plus_To_DataStream_en),
.proj_data_stream(PT_F1L5_Plus_To_DataStream),
.start(TPROJ_ToPlus_F3D5F4D5_F1_start),
.done(PT_F1L5_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L1L6F4") PT_L1L6F4_Plus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus_number),
.read_add_projin_disk_2(TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus_read_add),
.projin_disk_2(TPROJ_ToPlus_F1D5F2D5_F4_PT_L1L6F4_Plus),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_disk_8(6'b0),
.number_in_projin_disk_9(6'b0),
.number_in_projin_layer_1(6'b0),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(6'b0),
.number_in_projin_layer_5(6'b0),
.number_in_projin_layer_6(6'b0),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L1L6F4_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L1L6F4_Plus_From_DataStream),
.projout_disk_1(PT_L1L6F4_Plus_TPROJ_FromPlus_F4D5_F1F2),
.valid_disk_1(PT_L1L6F4_Plus_TPROJ_FromPlus_F4D5_F1F2_wr_en),
.valid_proj_data_stream(PT_L1L6F4_Plus_To_DataStream_en),
.proj_data_stream(PT_L1L6F4_Plus_To_DataStream),
.start(TPROJ_ToPlus_F1D5F2D5_F4_start),
.done(PT_L1L6F4_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L3F3F5") PT_L3F3F5_Minus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus_number),
.read_add_projin_disk_2(TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus_read_add),
.projin_disk_2(TPROJ_ToMinus_F1D5F2D5_F5_PT_L3F3F5_Minus),
.number_in_projin_disk_3(TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus_number),
.read_add_projin_disk_3(TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus_read_add),
.projin_disk_3(TPROJ_ToMinus_F3D5F4D5_F5_PT_L3F3F5_Minus),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus_number),
.read_add_projin_disk_7(TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus_read_add),
.projin_disk_7(TPROJ_ToMinus_F1D5F2D5_F3_PT_L3F3F5_Minus),
.number_in_projin_disk_8(6'b0),
.number_in_projin_disk_9(6'b0),
.number_in_projin_layer_1(6'b0),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(6'b0),
.number_in_projin_layer_5(6'b0),
.number_in_projin_layer_6(6'b0),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L3F3F5_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L3F3F5_Minus_From_DataStream),
.projout_disk_1(PT_L3F3F5_Minus_TPROJ_FromMinus_F3D5_F1F2),
.valid_disk_1(PT_L3F3F5_Minus_TPROJ_FromMinus_F3D5_F1F2_wr_en),
.projout_disk_3(PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F1F2),
.valid_disk_3(PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F1F2_wr_en),
.projout_disk_5(PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F3F4),
.valid_disk_5(PT_L3F3F5_Minus_TPROJ_FromMinus_F5D5_F3F4_wr_en),
.valid_proj_data_stream(PT_L3F3F5_Minus_To_DataStream_en),
.proj_data_stream(PT_L3F3F5_Minus_To_DataStream),
.start(TPROJ_ToMinus_F1D5F2D5_F5_start),
.done(PT_L3F3F5_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L2L4F2") PT_L2L4F2_Minus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus_number),
.read_add_projin_disk_2(TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus_read_add),
.projin_disk_2(TPROJ_ToMinus_F3D5F4D5_F2_PT_L2L4F2_Minus),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_disk_8(6'b0),
.number_in_projin_disk_9(6'b0),
.number_in_projin_layer_1(6'b0),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(6'b0),
.number_in_projin_layer_5(6'b0),
.number_in_projin_layer_6(6'b0),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L2L4F2_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L2L4F2_Minus_From_DataStream),
.projout_disk_1(PT_L2L4F2_Minus_TPROJ_FromMinus_F2D5_F3F4),
.valid_disk_1(PT_L2L4F2_Minus_TPROJ_FromMinus_F2D5_F3F4_wr_en),
.valid_proj_data_stream(PT_L2L4F2_Minus_To_DataStream_en),
.proj_data_stream(PT_L2L4F2_Minus_To_DataStream),
.start(TPROJ_ToMinus_F3D5F4D5_F2_start),
.done(PT_L2L4F2_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("F1L5") PT_F1L5_Minus(
.number_in_projin_disk_1(TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus_number),
.read_add_projin_disk_1(TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus_read_add),
.projin_disk_1(TPROJ_ToMinus_F3D5F4D5_F1_PT_F1L5_Minus),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_disk_8(6'b0),
.number_in_projin_disk_9(6'b0),
.number_in_projin_layer_1(6'b0),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(6'b0),
.number_in_projin_layer_5(6'b0),
.number_in_projin_layer_6(6'b0),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_F1L5_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_F1L5_Minus_From_DataStream),
.projout_disk_1(PT_F1L5_Minus_TPROJ_FromMinus_F1D5_F3F4),
.valid_disk_1(PT_F1L5_Minus_TPROJ_FromMinus_F1D5_F3F4_wr_en),
.valid_proj_data_stream(PT_F1L5_Minus_To_DataStream_en),
.proj_data_stream(PT_F1L5_Minus_To_DataStream),
.start(TPROJ_ToMinus_F3D5F4D5_F1_start),
.done(PT_F1L5_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L1L6F4") PT_L1L6F4_Minus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus_number),
.read_add_projin_disk_2(TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus_read_add),
.projin_disk_2(TPROJ_ToMinus_F1D5F2D5_F4_PT_L1L6F4_Minus),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_disk_8(6'b0),
.number_in_projin_disk_9(6'b0),
.number_in_projin_layer_1(6'b0),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(6'b0),
.number_in_projin_layer_5(6'b0),
.number_in_projin_layer_6(6'b0),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L1L6F4_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L1L6F4_Minus_From_DataStream),
.projout_disk_1(PT_L1L6F4_Minus_TPROJ_FromMinus_F4D5_F1F2),
.valid_disk_1(PT_L1L6F4_Minus_TPROJ_FromMinus_F4D5_F1F2_wr_en),
.valid_proj_data_stream(PT_L1L6F4_Minus_To_DataStream_en),
.proj_data_stream(PT_L1L6F4_Minus_To_DataStream),
.start(TPROJ_ToMinus_F1D5F2D5_F4_start),
.done(PT_L1L6F4_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  DR1_D5(
.stubin(IL1_D5_DR1_D5),
.stubout1(DR1_D5_SD1_F1D5),
.stubout2(DR1_D5_SD1_F2D5),
.stubout3(DR1_D5_SD1_F3D5),
.stubout4(DR1_D5_SD1_F4D5),
.stubout5(DR1_D5_SD1_F5D5),
.wr_en1(DR1_D5_SD1_F1D5_wr_en),
.wr_en2(DR1_D5_SD1_F2D5_wr_en),
.wr_en3(DR1_D5_SD1_F3D5_wr_en),
.wr_en4(DR1_D5_SD1_F4D5_wr_en),
.wr_en5(DR1_D5_SD1_F5D5_wr_en),
.start(IL1_D5_start),
.done(DR1_D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  DR2_D5(
.stubin(IL2_D5_DR2_D5),
.stubout1(DR2_D5_SD2_F1D5),
.stubout2(DR2_D5_SD2_F2D5),
.stubout3(DR2_D5_SD2_F3D5),
.stubout4(DR2_D5_SD2_F4D5),
.stubout5(DR2_D5_SD2_F5D5),
.wr_en1(DR2_D5_SD2_F1D5_wr_en),
.wr_en2(DR2_D5_SD2_F2D5_wr_en),
.wr_en3(DR2_D5_SD2_F3D5_wr_en),
.wr_en4(DR2_D5_SD2_F4D5_wr_en),
.wr_en5(DR2_D5_SD2_F5D5_wr_en),
.start(IL2_D5_start),
.done(DR2_D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  DR3_D5(
.stubin(IL3_D5_DR3_D5),
.stubout1(DR3_D5_SD3_F1D5),
.stubout2(DR3_D5_SD3_F2D5),
.stubout3(DR3_D5_SD3_F3D5),
.stubout4(DR3_D5_SD3_F4D5),
.stubout5(DR3_D5_SD3_F5D5),
.wr_en1(DR3_D5_SD3_F1D5_wr_en),
.wr_en2(DR3_D5_SD3_F2D5_wr_en),
.wr_en3(DR3_D5_SD3_F3D5_wr_en),
.wr_en4(DR3_D5_SD3_F4D5_wr_en),
.wr_en5(DR3_D5_SD3_F5D5_wr_en),
.start(IL3_D5_start),
.done(DR3_D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b1,1'b0) VMRD_F1D5(
.number_in_stubinLink1(SD1_F1D5_VMRD_F1D5_number),
.read_add_stubinLink1(SD1_F1D5_VMRD_F1D5_read_add),
.stubinLink1(SD1_F1D5_VMRD_F1D5),
.number_in_stubinLink2(SD2_F1D5_VMRD_F1D5_number),
.read_add_stubinLink2(SD2_F1D5_VMRD_F1D5_read_add),
.stubinLink2(SD2_F1D5_VMRD_F1D5),
.number_in_stubinLink3(SD3_F1D5_VMRD_F1D5_number),
.read_add_stubinLink3(SD3_F1D5_VMRD_F1D5_read_add),
.stubinLink3(SD3_F1D5_VMRD_F1D5),
.vmstuboutPHI1X1n1(VMRD_F1D5_VMS_F1D5PHI1X1n1),
.vmstuboutPHI1X1n2(VMRD_F1D5_VMS_F1D5PHI1X1n2),
.vmstuboutPHI1X1n3(VMRD_F1D5_VMS_F1D5PHI1X1n3),
.vmstuboutPHI2X1n1(VMRD_F1D5_VMS_F1D5PHI2X1n1),
.vmstuboutPHI2X1n2(VMRD_F1D5_VMS_F1D5PHI2X1n2),
.vmstuboutPHI2X1n3(VMRD_F1D5_VMS_F1D5PHI2X1n3),
.vmstuboutPHI2X1n4(VMRD_F1D5_VMS_F1D5PHI2X1n4),
.vmstuboutPHI2X1n5(VMRD_F1D5_VMS_F1D5PHI2X1n5),
.vmstuboutPHI3X1n1(VMRD_F1D5_VMS_F1D5PHI3X1n1),
.vmstuboutPHI3X1n2(VMRD_F1D5_VMS_F1D5PHI3X1n2),
.vmstuboutPHI3X1n3(VMRD_F1D5_VMS_F1D5PHI3X1n3),
.vmstuboutPHI3X1n4(VMRD_F1D5_VMS_F1D5PHI3X1n4),
.vmstuboutPHI3X1n5(VMRD_F1D5_VMS_F1D5PHI3X1n5),
.vmstuboutPHI4X1n1(VMRD_F1D5_VMS_F1D5PHI4X1n1),
.vmstuboutPHI4X1n2(VMRD_F1D5_VMS_F1D5PHI4X1n2),
.vmstuboutPHI4X1n3(VMRD_F1D5_VMS_F1D5PHI4X1n3),
.vmstuboutPHI1X2n1(VMRD_F1D5_VMS_F1D5PHI1X2n1),
.vmstuboutPHI1X2n2(VMRD_F1D5_VMS_F1D5PHI1X2n2),
.vmstuboutPHI2X2n1(VMRD_F1D5_VMS_F1D5PHI2X2n1),
.vmstuboutPHI2X2n2(VMRD_F1D5_VMS_F1D5PHI2X2n2),
.vmstuboutPHI2X2n3(VMRD_F1D5_VMS_F1D5PHI2X2n3),
.vmstuboutPHI3X2n1(VMRD_F1D5_VMS_F1D5PHI3X2n1),
.vmstuboutPHI3X2n2(VMRD_F1D5_VMS_F1D5PHI3X2n2),
.vmstuboutPHI3X2n3(VMRD_F1D5_VMS_F1D5PHI3X2n3),
.vmstuboutPHI4X2n1(VMRD_F1D5_VMS_F1D5PHI4X2n1),
.vmstuboutPHI4X2n2(VMRD_F1D5_VMS_F1D5PHI4X2n2),
.allstuboutn1(VMRD_F1D5_AS_F1D5n1),
.allstuboutn2(VMRD_F1D5_AS_F1D5n2),
.vmstuboutPHI1X1n1_wr_en(VMRD_F1D5_VMS_F1D5PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMRD_F1D5_VMS_F1D5PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMRD_F1D5_VMS_F1D5PHI1X1n3_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMRD_F1D5_VMS_F1D5PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMRD_F1D5_VMS_F1D5PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMRD_F1D5_VMS_F1D5PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMRD_F1D5_VMS_F1D5PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMRD_F1D5_VMS_F1D5PHI2X1n5_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMRD_F1D5_VMS_F1D5PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMRD_F1D5_VMS_F1D5PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMRD_F1D5_VMS_F1D5PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMRD_F1D5_VMS_F1D5PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMRD_F1D5_VMS_F1D5PHI3X1n5_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMRD_F1D5_VMS_F1D5PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMRD_F1D5_VMS_F1D5PHI4X1n2_wr_en),
.vmstuboutPHI4X1n3_wr_en(VMRD_F1D5_VMS_F1D5PHI4X1n3_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMRD_F1D5_VMS_F1D5PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMRD_F1D5_VMS_F1D5PHI1X2n2_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMRD_F1D5_VMS_F1D5PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMRD_F1D5_VMS_F1D5PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMRD_F1D5_VMS_F1D5PHI2X2n3_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMRD_F1D5_VMS_F1D5PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMRD_F1D5_VMS_F1D5PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMRD_F1D5_VMS_F1D5PHI3X2n3_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMRD_F1D5_VMS_F1D5PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMRD_F1D5_VMS_F1D5PHI4X2n2_wr_en),
.valid_data1(VMRD_F1D5_AS_F1D5n1_wr_en),
.valid_data2(VMRD_F1D5_AS_F1D5n2_wr_en),
.start(SD1_F1D5_start),
.done(VMRD_F1D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b0,1'b0) VMRD_F2D5(
.number_in_stubinLink1(SD1_F2D5_VMRD_F2D5_number),
.read_add_stubinLink1(SD1_F2D5_VMRD_F2D5_read_add),
.stubinLink1(SD1_F2D5_VMRD_F2D5),
.number_in_stubinLink2(SD2_F2D5_VMRD_F2D5_number),
.read_add_stubinLink2(SD2_F2D5_VMRD_F2D5_read_add),
.stubinLink2(SD2_F2D5_VMRD_F2D5),
.number_in_stubinLink3(SD3_F2D5_VMRD_F2D5_number),
.read_add_stubinLink3(SD3_F2D5_VMRD_F2D5_read_add),
.stubinLink3(SD3_F2D5_VMRD_F2D5),
.vmstuboutPHI1X1n1(VMRD_F2D5_VMS_F2D5PHI1X1n1),
.vmstuboutPHI1X1n2(VMRD_F2D5_VMS_F2D5PHI1X1n2),
.vmstuboutPHI1X1n3(VMRD_F2D5_VMS_F2D5PHI1X1n3),
.vmstuboutPHI2X1n1(VMRD_F2D5_VMS_F2D5PHI2X1n1),
.vmstuboutPHI2X1n2(VMRD_F2D5_VMS_F2D5PHI2X1n2),
.vmstuboutPHI2X1n3(VMRD_F2D5_VMS_F2D5PHI2X1n3),
.vmstuboutPHI3X1n1(VMRD_F2D5_VMS_F2D5PHI3X1n1),
.vmstuboutPHI3X1n2(VMRD_F2D5_VMS_F2D5PHI3X1n2),
.vmstuboutPHI3X1n3(VMRD_F2D5_VMS_F2D5PHI3X1n3),
.vmstuboutPHI1X2n1(VMRD_F2D5_VMS_F2D5PHI1X2n1),
.vmstuboutPHI1X2n2(VMRD_F2D5_VMS_F2D5PHI1X2n2),
.vmstuboutPHI1X2n3(VMRD_F2D5_VMS_F2D5PHI1X2n3),
.vmstuboutPHI1X2n4(VMRD_F2D5_VMS_F2D5PHI1X2n4),
.vmstuboutPHI1X2n5(VMRD_F2D5_VMS_F2D5PHI1X2n5),
.vmstuboutPHI2X2n1(VMRD_F2D5_VMS_F2D5PHI2X2n1),
.vmstuboutPHI2X2n2(VMRD_F2D5_VMS_F2D5PHI2X2n2),
.vmstuboutPHI2X2n3(VMRD_F2D5_VMS_F2D5PHI2X2n3),
.vmstuboutPHI2X2n4(VMRD_F2D5_VMS_F2D5PHI2X2n4),
.vmstuboutPHI2X2n5(VMRD_F2D5_VMS_F2D5PHI2X2n5),
.vmstuboutPHI3X2n1(VMRD_F2D5_VMS_F2D5PHI3X2n1),
.vmstuboutPHI3X2n2(VMRD_F2D5_VMS_F2D5PHI3X2n2),
.vmstuboutPHI3X2n3(VMRD_F2D5_VMS_F2D5PHI3X2n3),
.vmstuboutPHI3X2n4(VMRD_F2D5_VMS_F2D5PHI3X2n4),
.vmstuboutPHI3X2n5(VMRD_F2D5_VMS_F2D5PHI3X2n5),
.allstuboutn1(VMRD_F2D5_AS_F2D5n1),
.allstuboutn2(VMRD_F2D5_AS_F2D5n2),
.vmstuboutPHI1X1n1_wr_en(VMRD_F2D5_VMS_F2D5PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMRD_F2D5_VMS_F2D5PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMRD_F2D5_VMS_F2D5PHI1X1n3_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMRD_F2D5_VMS_F2D5PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMRD_F2D5_VMS_F2D5PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMRD_F2D5_VMS_F2D5PHI2X1n3_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMRD_F2D5_VMS_F2D5PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMRD_F2D5_VMS_F2D5PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMRD_F2D5_VMS_F2D5PHI3X1n3_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMRD_F2D5_VMS_F2D5PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMRD_F2D5_VMS_F2D5PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMRD_F2D5_VMS_F2D5PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMRD_F2D5_VMS_F2D5PHI1X2n4_wr_en),
.vmstuboutPHI1X2n5_wr_en(VMRD_F2D5_VMS_F2D5PHI1X2n5_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMRD_F2D5_VMS_F2D5PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMRD_F2D5_VMS_F2D5PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMRD_F2D5_VMS_F2D5PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMRD_F2D5_VMS_F2D5PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMRD_F2D5_VMS_F2D5PHI2X2n5_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMRD_F2D5_VMS_F2D5PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMRD_F2D5_VMS_F2D5PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMRD_F2D5_VMS_F2D5PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMRD_F2D5_VMS_F2D5PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMRD_F2D5_VMS_F2D5PHI3X2n5_wr_en),
.valid_data1(VMRD_F2D5_AS_F2D5n1_wr_en),
.valid_data2(VMRD_F2D5_AS_F2D5n2_wr_en),
.start(SD1_F2D5_start),
.done(VMRD_F2D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b1,1'b0) VMRD_F3D5(
.number_in_stubinLink1(SD1_F3D5_VMRD_F3D5_number),
.read_add_stubinLink1(SD1_F3D5_VMRD_F3D5_read_add),
.stubinLink1(SD1_F3D5_VMRD_F3D5),
.number_in_stubinLink2(SD2_F3D5_VMRD_F3D5_number),
.read_add_stubinLink2(SD2_F3D5_VMRD_F3D5_read_add),
.stubinLink2(SD2_F3D5_VMRD_F3D5),
.number_in_stubinLink3(SD3_F3D5_VMRD_F3D5_number),
.read_add_stubinLink3(SD3_F3D5_VMRD_F3D5_read_add),
.stubinLink3(SD3_F3D5_VMRD_F3D5),
.vmstuboutPHI1X1n1(VMRD_F3D5_VMS_F3D5PHI1X1n1),
.vmstuboutPHI1X1n2(VMRD_F3D5_VMS_F3D5PHI1X1n2),
.vmstuboutPHI1X1n3(VMRD_F3D5_VMS_F3D5PHI1X1n3),
.vmstuboutPHI2X1n1(VMRD_F3D5_VMS_F3D5PHI2X1n1),
.vmstuboutPHI2X1n2(VMRD_F3D5_VMS_F3D5PHI2X1n2),
.vmstuboutPHI2X1n3(VMRD_F3D5_VMS_F3D5PHI2X1n3),
.vmstuboutPHI2X1n4(VMRD_F3D5_VMS_F3D5PHI2X1n4),
.vmstuboutPHI2X1n5(VMRD_F3D5_VMS_F3D5PHI2X1n5),
.vmstuboutPHI3X1n1(VMRD_F3D5_VMS_F3D5PHI3X1n1),
.vmstuboutPHI3X1n2(VMRD_F3D5_VMS_F3D5PHI3X1n2),
.vmstuboutPHI3X1n3(VMRD_F3D5_VMS_F3D5PHI3X1n3),
.vmstuboutPHI3X1n4(VMRD_F3D5_VMS_F3D5PHI3X1n4),
.vmstuboutPHI3X1n5(VMRD_F3D5_VMS_F3D5PHI3X1n5),
.vmstuboutPHI4X1n1(VMRD_F3D5_VMS_F3D5PHI4X1n1),
.vmstuboutPHI4X1n2(VMRD_F3D5_VMS_F3D5PHI4X1n2),
.vmstuboutPHI4X1n3(VMRD_F3D5_VMS_F3D5PHI4X1n3),
.vmstuboutPHI1X2n1(VMRD_F3D5_VMS_F3D5PHI1X2n1),
.vmstuboutPHI1X2n2(VMRD_F3D5_VMS_F3D5PHI1X2n2),
.vmstuboutPHI2X2n1(VMRD_F3D5_VMS_F3D5PHI2X2n1),
.vmstuboutPHI2X2n2(VMRD_F3D5_VMS_F3D5PHI2X2n2),
.vmstuboutPHI2X2n3(VMRD_F3D5_VMS_F3D5PHI2X2n3),
.vmstuboutPHI3X2n1(VMRD_F3D5_VMS_F3D5PHI3X2n1),
.vmstuboutPHI3X2n2(VMRD_F3D5_VMS_F3D5PHI3X2n2),
.vmstuboutPHI3X2n3(VMRD_F3D5_VMS_F3D5PHI3X2n3),
.vmstuboutPHI4X2n1(VMRD_F3D5_VMS_F3D5PHI4X2n1),
.vmstuboutPHI4X2n2(VMRD_F3D5_VMS_F3D5PHI4X2n2),
.allstuboutn1(VMRD_F3D5_AS_F3D5n1),
.allstuboutn2(VMRD_F3D5_AS_F3D5n2),
.vmstuboutPHI1X1n1_wr_en(VMRD_F3D5_VMS_F3D5PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMRD_F3D5_VMS_F3D5PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMRD_F3D5_VMS_F3D5PHI1X1n3_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMRD_F3D5_VMS_F3D5PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMRD_F3D5_VMS_F3D5PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMRD_F3D5_VMS_F3D5PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMRD_F3D5_VMS_F3D5PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMRD_F3D5_VMS_F3D5PHI2X1n5_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMRD_F3D5_VMS_F3D5PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMRD_F3D5_VMS_F3D5PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMRD_F3D5_VMS_F3D5PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMRD_F3D5_VMS_F3D5PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMRD_F3D5_VMS_F3D5PHI3X1n5_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMRD_F3D5_VMS_F3D5PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMRD_F3D5_VMS_F3D5PHI4X1n2_wr_en),
.vmstuboutPHI4X1n3_wr_en(VMRD_F3D5_VMS_F3D5PHI4X1n3_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMRD_F3D5_VMS_F3D5PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMRD_F3D5_VMS_F3D5PHI1X2n2_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMRD_F3D5_VMS_F3D5PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMRD_F3D5_VMS_F3D5PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMRD_F3D5_VMS_F3D5PHI2X2n3_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMRD_F3D5_VMS_F3D5PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMRD_F3D5_VMS_F3D5PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMRD_F3D5_VMS_F3D5PHI3X2n3_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMRD_F3D5_VMS_F3D5PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMRD_F3D5_VMS_F3D5PHI4X2n2_wr_en),
.valid_data1(VMRD_F3D5_AS_F3D5n1_wr_en),
.valid_data2(VMRD_F3D5_AS_F3D5n2_wr_en),
.start(SD1_F3D5_start),
.done(VMRD_F3D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b0,1'b0) VMRD_F4D5(
.number_in_stubinLink1(SD1_F4D5_VMRD_F4D5_number),
.read_add_stubinLink1(SD1_F4D5_VMRD_F4D5_read_add),
.stubinLink1(SD1_F4D5_VMRD_F4D5),
.number_in_stubinLink2(SD2_F4D5_VMRD_F4D5_number),
.read_add_stubinLink2(SD2_F4D5_VMRD_F4D5_read_add),
.stubinLink2(SD2_F4D5_VMRD_F4D5),
.number_in_stubinLink3(SD3_F4D5_VMRD_F4D5_number),
.read_add_stubinLink3(SD3_F4D5_VMRD_F4D5_read_add),
.stubinLink3(SD3_F4D5_VMRD_F4D5),
.vmstuboutPHI1X1n1(VMRD_F4D5_VMS_F4D5PHI1X1n1),
.vmstuboutPHI1X1n2(VMRD_F4D5_VMS_F4D5PHI1X1n2),
.vmstuboutPHI1X1n3(VMRD_F4D5_VMS_F4D5PHI1X1n3),
.vmstuboutPHI2X1n1(VMRD_F4D5_VMS_F4D5PHI2X1n1),
.vmstuboutPHI2X1n2(VMRD_F4D5_VMS_F4D5PHI2X1n2),
.vmstuboutPHI2X1n3(VMRD_F4D5_VMS_F4D5PHI2X1n3),
.vmstuboutPHI3X1n1(VMRD_F4D5_VMS_F4D5PHI3X1n1),
.vmstuboutPHI3X1n2(VMRD_F4D5_VMS_F4D5PHI3X1n2),
.vmstuboutPHI3X1n3(VMRD_F4D5_VMS_F4D5PHI3X1n3),
.vmstuboutPHI1X2n1(VMRD_F4D5_VMS_F4D5PHI1X2n1),
.vmstuboutPHI1X2n2(VMRD_F4D5_VMS_F4D5PHI1X2n2),
.vmstuboutPHI1X2n3(VMRD_F4D5_VMS_F4D5PHI1X2n3),
.vmstuboutPHI1X2n4(VMRD_F4D5_VMS_F4D5PHI1X2n4),
.vmstuboutPHI1X2n5(VMRD_F4D5_VMS_F4D5PHI1X2n5),
.vmstuboutPHI2X2n1(VMRD_F4D5_VMS_F4D5PHI2X2n1),
.vmstuboutPHI2X2n2(VMRD_F4D5_VMS_F4D5PHI2X2n2),
.vmstuboutPHI2X2n3(VMRD_F4D5_VMS_F4D5PHI2X2n3),
.vmstuboutPHI2X2n4(VMRD_F4D5_VMS_F4D5PHI2X2n4),
.vmstuboutPHI2X2n5(VMRD_F4D5_VMS_F4D5PHI2X2n5),
.vmstuboutPHI3X2n1(VMRD_F4D5_VMS_F4D5PHI3X2n1),
.vmstuboutPHI3X2n2(VMRD_F4D5_VMS_F4D5PHI3X2n2),
.vmstuboutPHI3X2n3(VMRD_F4D5_VMS_F4D5PHI3X2n3),
.vmstuboutPHI3X2n4(VMRD_F4D5_VMS_F4D5PHI3X2n4),
.vmstuboutPHI3X2n5(VMRD_F4D5_VMS_F4D5PHI3X2n5),
.allstuboutn1(VMRD_F4D5_AS_F4D5n1),
.allstuboutn2(VMRD_F4D5_AS_F4D5n2),
.vmstuboutPHI1X1n1_wr_en(VMRD_F4D5_VMS_F4D5PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMRD_F4D5_VMS_F4D5PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMRD_F4D5_VMS_F4D5PHI1X1n3_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMRD_F4D5_VMS_F4D5PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMRD_F4D5_VMS_F4D5PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMRD_F4D5_VMS_F4D5PHI2X1n3_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMRD_F4D5_VMS_F4D5PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMRD_F4D5_VMS_F4D5PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMRD_F4D5_VMS_F4D5PHI3X1n3_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMRD_F4D5_VMS_F4D5PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMRD_F4D5_VMS_F4D5PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMRD_F4D5_VMS_F4D5PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMRD_F4D5_VMS_F4D5PHI1X2n4_wr_en),
.vmstuboutPHI1X2n5_wr_en(VMRD_F4D5_VMS_F4D5PHI1X2n5_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMRD_F4D5_VMS_F4D5PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMRD_F4D5_VMS_F4D5PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMRD_F4D5_VMS_F4D5PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMRD_F4D5_VMS_F4D5PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMRD_F4D5_VMS_F4D5PHI2X2n5_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMRD_F4D5_VMS_F4D5PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMRD_F4D5_VMS_F4D5PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMRD_F4D5_VMS_F4D5PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMRD_F4D5_VMS_F4D5PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMRD_F4D5_VMS_F4D5PHI3X2n5_wr_en),
.valid_data1(VMRD_F4D5_AS_F4D5n1_wr_en),
.valid_data2(VMRD_F4D5_AS_F4D5n2_wr_en),
.start(SD1_F4D5_start),
.done(VMRD_F4D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b1,1'b0) VMRD_F5D5(
.number_in_stubinLink1(SD1_F5D5_VMRD_F5D5_number),
.read_add_stubinLink1(SD1_F5D5_VMRD_F5D5_read_add),
.stubinLink1(SD1_F5D5_VMRD_F5D5),
.number_in_stubinLink2(SD2_F5D5_VMRD_F5D5_number),
.read_add_stubinLink2(SD2_F5D5_VMRD_F5D5_read_add),
.stubinLink2(SD2_F5D5_VMRD_F5D5),
.number_in_stubinLink3(SD3_F5D5_VMRD_F5D5_number),
.read_add_stubinLink3(SD3_F5D5_VMRD_F5D5_read_add),
.stubinLink3(SD3_F5D5_VMRD_F5D5),
.vmstuboutPHI1X1n1(VMRD_F5D5_VMS_F5D5PHI1X1n1),
.vmstuboutPHI1X1n2(VMRD_F5D5_VMS_F5D5PHI1X1n2),
.vmstuboutPHI1X2n1(VMRD_F5D5_VMS_F5D5PHI1X2n1),
.vmstuboutPHI1X2n2(VMRD_F5D5_VMS_F5D5PHI1X2n2),
.vmstuboutPHI2X1n1(VMRD_F5D5_VMS_F5D5PHI2X1n1),
.vmstuboutPHI2X1n2(VMRD_F5D5_VMS_F5D5PHI2X1n2),
.vmstuboutPHI2X2n1(VMRD_F5D5_VMS_F5D5PHI2X2n1),
.vmstuboutPHI2X2n2(VMRD_F5D5_VMS_F5D5PHI2X2n2),
.vmstuboutPHI3X1n1(VMRD_F5D5_VMS_F5D5PHI3X1n1),
.vmstuboutPHI3X1n2(VMRD_F5D5_VMS_F5D5PHI3X1n2),
.vmstuboutPHI3X2n1(VMRD_F5D5_VMS_F5D5PHI3X2n1),
.vmstuboutPHI3X2n2(VMRD_F5D5_VMS_F5D5PHI3X2n2),
.vmstuboutPHI4X1n1(VMRD_F5D5_VMS_F5D5PHI4X1n1),
.vmstuboutPHI4X1n2(VMRD_F5D5_VMS_F5D5PHI4X1n2),
.vmstuboutPHI4X2n1(VMRD_F5D5_VMS_F5D5PHI4X2n1),
.vmstuboutPHI4X2n2(VMRD_F5D5_VMS_F5D5PHI4X2n2),
.allstuboutn1(VMRD_F5D5_AS_F5D5n1),
.allstuboutn2(VMRD_F5D5_AS_F5D5n2),
.vmstuboutPHI1X1n1_wr_en(VMRD_F5D5_VMS_F5D5PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMRD_F5D5_VMS_F5D5PHI1X1n2_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMRD_F5D5_VMS_F5D5PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMRD_F5D5_VMS_F5D5PHI1X2n2_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMRD_F5D5_VMS_F5D5PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMRD_F5D5_VMS_F5D5PHI2X1n2_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMRD_F5D5_VMS_F5D5PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMRD_F5D5_VMS_F5D5PHI2X2n2_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMRD_F5D5_VMS_F5D5PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMRD_F5D5_VMS_F5D5PHI3X1n2_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMRD_F5D5_VMS_F5D5PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMRD_F5D5_VMS_F5D5PHI3X2n2_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMRD_F5D5_VMS_F5D5PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMRD_F5D5_VMS_F5D5PHI4X1n2_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMRD_F5D5_VMS_F5D5PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMRD_F5D5_VMS_F5D5PHI4X2n2_wr_en),
.valid_data1(VMRD_F5D5_AS_F5D5n1_wr_en),
.valid_data2(VMRD_F5D5_AS_F5D5n2_wr_en),
.start(SD1_F5D5_start),
.done(VMRD_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI1X1_F2D5PHI1X1_phi.txt","TETable_TE_F1D5PHI1X1_F2D5PHI1X1_z.txt",1'b0) TE_F1D5PHI1X1_F2D5PHI1X1(
.number_in_innervmstubin(VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_number),
.read_add_innervmstubin(VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_read_add),
.innervmstubin(VMS_F1D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1),
.number_in_outervmstubin(VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_number),
.read_add_outervmstubin(VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1_read_add),
.outervmstubin(VMS_F2D5PHI1X1n1_TE_F1D5PHI1X1_F2D5PHI1X1),
.stubpairout(TE_F1D5PHI1X1_F2D5PHI1X1_SP_F1D5PHI1X1_F2D5PHI1X1),
.valid_data(TE_F1D5PHI1X1_F2D5PHI1X1_SP_F1D5PHI1X1_F2D5PHI1X1_wr_en),
.start(VMS_F1D5PHI1X1n1_start),
.done(TE_F1D5PHI1X1_F2D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI2X1_F2D5PHI1X1_phi.txt","TETable_TE_F1D5PHI2X1_F2D5PHI1X1_z.txt",1'b0) TE_F1D5PHI2X1_F2D5PHI1X1(
.number_in_outervmstubin(VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1_number),
.read_add_outervmstubin(VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1_read_add),
.outervmstubin(VMS_F2D5PHI1X1n2_TE_F1D5PHI2X1_F2D5PHI1X1),
.number_in_innervmstubin(VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1_number),
.read_add_innervmstubin(VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1_read_add),
.innervmstubin(VMS_F1D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI1X1),
.stubpairout(TE_F1D5PHI2X1_F2D5PHI1X1_SP_F1D5PHI2X1_F2D5PHI1X1),
.valid_data(TE_F1D5PHI2X1_F2D5PHI1X1_SP_F1D5PHI2X1_F2D5PHI1X1_wr_en),
.start(VMS_F2D5PHI1X1n2_start),
.done(TE_F1D5PHI2X1_F2D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI2X1_F2D5PHI2X1_phi.txt","TETable_TE_F1D5PHI2X1_F2D5PHI2X1_z.txt",1'b0) TE_F1D5PHI2X1_F2D5PHI2X1(
.number_in_innervmstubin(VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1_number),
.read_add_innervmstubin(VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1_read_add),
.innervmstubin(VMS_F1D5PHI2X1n2_TE_F1D5PHI2X1_F2D5PHI2X1),
.number_in_outervmstubin(VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1_number),
.read_add_outervmstubin(VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1_read_add),
.outervmstubin(VMS_F2D5PHI2X1n1_TE_F1D5PHI2X1_F2D5PHI2X1),
.stubpairout(TE_F1D5PHI2X1_F2D5PHI2X1_SP_F1D5PHI2X1_F2D5PHI2X1),
.valid_data(TE_F1D5PHI2X1_F2D5PHI2X1_SP_F1D5PHI2X1_F2D5PHI2X1_wr_en),
.start(VMS_F1D5PHI2X1n2_start),
.done(TE_F1D5PHI2X1_F2D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI3X1_F2D5PHI2X1_phi.txt","TETable_TE_F1D5PHI3X1_F2D5PHI2X1_z.txt",1'b0) TE_F1D5PHI3X1_F2D5PHI2X1(
.number_in_outervmstubin(VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1_number),
.read_add_outervmstubin(VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1_read_add),
.outervmstubin(VMS_F2D5PHI2X1n2_TE_F1D5PHI3X1_F2D5PHI2X1),
.number_in_innervmstubin(VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1_number),
.read_add_innervmstubin(VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1_read_add),
.innervmstubin(VMS_F1D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI2X1),
.stubpairout(TE_F1D5PHI3X1_F2D5PHI2X1_SP_F1D5PHI3X1_F2D5PHI2X1),
.valid_data(TE_F1D5PHI3X1_F2D5PHI2X1_SP_F1D5PHI3X1_F2D5PHI2X1_wr_en),
.start(VMS_F2D5PHI2X1n2_start),
.done(TE_F1D5PHI3X1_F2D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI3X1_F2D5PHI3X1_phi.txt","TETable_TE_F1D5PHI3X1_F2D5PHI3X1_z.txt",1'b0) TE_F1D5PHI3X1_F2D5PHI3X1(
.number_in_innervmstubin(VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1_number),
.read_add_innervmstubin(VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1_read_add),
.innervmstubin(VMS_F1D5PHI3X1n2_TE_F1D5PHI3X1_F2D5PHI3X1),
.number_in_outervmstubin(VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1_number),
.read_add_outervmstubin(VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1_read_add),
.outervmstubin(VMS_F2D5PHI3X1n1_TE_F1D5PHI3X1_F2D5PHI3X1),
.stubpairout(TE_F1D5PHI3X1_F2D5PHI3X1_SP_F1D5PHI3X1_F2D5PHI3X1),
.valid_data(TE_F1D5PHI3X1_F2D5PHI3X1_SP_F1D5PHI3X1_F2D5PHI3X1_wr_en),
.start(VMS_F1D5PHI3X1n2_start),
.done(TE_F1D5PHI3X1_F2D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI4X1_F2D5PHI3X1_phi.txt","TETable_TE_F1D5PHI4X1_F2D5PHI3X1_z.txt",1'b0) TE_F1D5PHI4X1_F2D5PHI3X1(
.number_in_outervmstubin(VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1_number),
.read_add_outervmstubin(VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1_read_add),
.outervmstubin(VMS_F2D5PHI3X1n2_TE_F1D5PHI4X1_F2D5PHI3X1),
.number_in_innervmstubin(VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1_number),
.read_add_innervmstubin(VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1_read_add),
.innervmstubin(VMS_F1D5PHI4X1n1_TE_F1D5PHI4X1_F2D5PHI3X1),
.stubpairout(TE_F1D5PHI4X1_F2D5PHI3X1_SP_F1D5PHI4X1_F2D5PHI3X1),
.valid_data(TE_F1D5PHI4X1_F2D5PHI3X1_SP_F1D5PHI4X1_F2D5PHI3X1_wr_en),
.start(VMS_F2D5PHI3X1n2_start),
.done(TE_F1D5PHI4X1_F2D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI1X1_F2D5PHI1X2_phi.txt","TETable_TE_F1D5PHI1X1_F2D5PHI1X2_z.txt",1'b0) TE_F1D5PHI1X1_F2D5PHI1X2(
.number_in_innervmstubin(VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2_number),
.read_add_innervmstubin(VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2_read_add),
.innervmstubin(VMS_F1D5PHI1X1n2_TE_F1D5PHI1X1_F2D5PHI1X2),
.number_in_outervmstubin(VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2_number),
.read_add_outervmstubin(VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2_read_add),
.outervmstubin(VMS_F2D5PHI1X2n1_TE_F1D5PHI1X1_F2D5PHI1X2),
.stubpairout(TE_F1D5PHI1X1_F2D5PHI1X2_SP_F1D5PHI1X1_F2D5PHI1X2),
.valid_data(TE_F1D5PHI1X1_F2D5PHI1X2_SP_F1D5PHI1X1_F2D5PHI1X2_wr_en),
.start(VMS_F1D5PHI1X1n2_start),
.done(TE_F1D5PHI1X1_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI2X1_F2D5PHI1X2_phi.txt","TETable_TE_F1D5PHI2X1_F2D5PHI1X2_z.txt",1'b0) TE_F1D5PHI2X1_F2D5PHI1X2(
.number_in_innervmstubin(VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2_number),
.read_add_innervmstubin(VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2_read_add),
.innervmstubin(VMS_F1D5PHI2X1n3_TE_F1D5PHI2X1_F2D5PHI1X2),
.number_in_outervmstubin(VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2_number),
.read_add_outervmstubin(VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2_read_add),
.outervmstubin(VMS_F2D5PHI1X2n2_TE_F1D5PHI2X1_F2D5PHI1X2),
.stubpairout(TE_F1D5PHI2X1_F2D5PHI1X2_SP_F1D5PHI2X1_F2D5PHI1X2),
.valid_data(TE_F1D5PHI2X1_F2D5PHI1X2_SP_F1D5PHI2X1_F2D5PHI1X2_wr_en),
.start(VMS_F1D5PHI2X1n3_start),
.done(TE_F1D5PHI2X1_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI2X1_F2D5PHI2X2_phi.txt","TETable_TE_F1D5PHI2X1_F2D5PHI2X2_z.txt",1'b0) TE_F1D5PHI2X1_F2D5PHI2X2(
.number_in_innervmstubin(VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2_number),
.read_add_innervmstubin(VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2_read_add),
.innervmstubin(VMS_F1D5PHI2X1n4_TE_F1D5PHI2X1_F2D5PHI2X2),
.number_in_outervmstubin(VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2_number),
.read_add_outervmstubin(VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2_read_add),
.outervmstubin(VMS_F2D5PHI2X2n1_TE_F1D5PHI2X1_F2D5PHI2X2),
.stubpairout(TE_F1D5PHI2X1_F2D5PHI2X2_SP_F1D5PHI2X1_F2D5PHI2X2),
.valid_data(TE_F1D5PHI2X1_F2D5PHI2X2_SP_F1D5PHI2X1_F2D5PHI2X2_wr_en),
.start(VMS_F1D5PHI2X1n4_start),
.done(TE_F1D5PHI2X1_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI3X1_F2D5PHI2X2_phi.txt","TETable_TE_F1D5PHI3X1_F2D5PHI2X2_z.txt",1'b0) TE_F1D5PHI3X1_F2D5PHI2X2(
.number_in_innervmstubin(VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2_number),
.read_add_innervmstubin(VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2_read_add),
.innervmstubin(VMS_F1D5PHI3X1n3_TE_F1D5PHI3X1_F2D5PHI2X2),
.number_in_outervmstubin(VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2_number),
.read_add_outervmstubin(VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2_read_add),
.outervmstubin(VMS_F2D5PHI2X2n2_TE_F1D5PHI3X1_F2D5PHI2X2),
.stubpairout(TE_F1D5PHI3X1_F2D5PHI2X2_SP_F1D5PHI3X1_F2D5PHI2X2),
.valid_data(TE_F1D5PHI3X1_F2D5PHI2X2_SP_F1D5PHI3X1_F2D5PHI2X2_wr_en),
.start(VMS_F1D5PHI3X1n3_start),
.done(TE_F1D5PHI3X1_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI3X1_F2D5PHI3X2_phi.txt","TETable_TE_F1D5PHI3X1_F2D5PHI3X2_z.txt",1'b0) TE_F1D5PHI3X1_F2D5PHI3X2(
.number_in_innervmstubin(VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2_number),
.read_add_innervmstubin(VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2_read_add),
.innervmstubin(VMS_F1D5PHI3X1n4_TE_F1D5PHI3X1_F2D5PHI3X2),
.number_in_outervmstubin(VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2_number),
.read_add_outervmstubin(VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2_read_add),
.outervmstubin(VMS_F2D5PHI3X2n1_TE_F1D5PHI3X1_F2D5PHI3X2),
.stubpairout(TE_F1D5PHI3X1_F2D5PHI3X2_SP_F1D5PHI3X1_F2D5PHI3X2),
.valid_data(TE_F1D5PHI3X1_F2D5PHI3X2_SP_F1D5PHI3X1_F2D5PHI3X2_wr_en),
.start(VMS_F1D5PHI3X1n4_start),
.done(TE_F1D5PHI3X1_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI4X1_F2D5PHI3X2_phi.txt","TETable_TE_F1D5PHI4X1_F2D5PHI3X2_z.txt",1'b0) TE_F1D5PHI4X1_F2D5PHI3X2(
.number_in_innervmstubin(VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2_number),
.read_add_innervmstubin(VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2_read_add),
.innervmstubin(VMS_F1D5PHI4X1n2_TE_F1D5PHI4X1_F2D5PHI3X2),
.number_in_outervmstubin(VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2_number),
.read_add_outervmstubin(VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2_read_add),
.outervmstubin(VMS_F2D5PHI3X2n2_TE_F1D5PHI4X1_F2D5PHI3X2),
.stubpairout(TE_F1D5PHI4X1_F2D5PHI3X2_SP_F1D5PHI4X1_F2D5PHI3X2),
.valid_data(TE_F1D5PHI4X1_F2D5PHI3X2_SP_F1D5PHI4X1_F2D5PHI3X2_wr_en),
.start(VMS_F1D5PHI4X1n2_start),
.done(TE_F1D5PHI4X1_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI1X2_F2D5PHI1X2_phi.txt","TETable_TE_F1D5PHI1X2_F2D5PHI1X2_z.txt",1'b0) TE_F1D5PHI1X2_F2D5PHI1X2(
.number_in_outervmstubin(VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2_number),
.read_add_outervmstubin(VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2_read_add),
.outervmstubin(VMS_F2D5PHI1X2n3_TE_F1D5PHI1X2_F2D5PHI1X2),
.number_in_innervmstubin(VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2_number),
.read_add_innervmstubin(VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2_read_add),
.innervmstubin(VMS_F1D5PHI1X2n1_TE_F1D5PHI1X2_F2D5PHI1X2),
.stubpairout(TE_F1D5PHI1X2_F2D5PHI1X2_SP_F1D5PHI1X2_F2D5PHI1X2),
.valid_data(TE_F1D5PHI1X2_F2D5PHI1X2_SP_F1D5PHI1X2_F2D5PHI1X2_wr_en),
.start(VMS_F2D5PHI1X2n3_start),
.done(TE_F1D5PHI1X2_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI2X2_F2D5PHI1X2_phi.txt","TETable_TE_F1D5PHI2X2_F2D5PHI1X2_z.txt",1'b0) TE_F1D5PHI2X2_F2D5PHI1X2(
.number_in_outervmstubin(VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2_number),
.read_add_outervmstubin(VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2_read_add),
.outervmstubin(VMS_F2D5PHI1X2n4_TE_F1D5PHI2X2_F2D5PHI1X2),
.number_in_innervmstubin(VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2_number),
.read_add_innervmstubin(VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2_read_add),
.innervmstubin(VMS_F1D5PHI2X2n1_TE_F1D5PHI2X2_F2D5PHI1X2),
.stubpairout(TE_F1D5PHI2X2_F2D5PHI1X2_SP_F1D5PHI2X2_F2D5PHI1X2),
.valid_data(TE_F1D5PHI2X2_F2D5PHI1X2_SP_F1D5PHI2X2_F2D5PHI1X2_wr_en),
.start(VMS_F2D5PHI1X2n4_start),
.done(TE_F1D5PHI2X2_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI2X2_F2D5PHI2X2_phi.txt","TETable_TE_F1D5PHI2X2_F2D5PHI2X2_z.txt",1'b0) TE_F1D5PHI2X2_F2D5PHI2X2(
.number_in_outervmstubin(VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2_number),
.read_add_outervmstubin(VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2_read_add),
.outervmstubin(VMS_F2D5PHI2X2n3_TE_F1D5PHI2X2_F2D5PHI2X2),
.number_in_innervmstubin(VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2_number),
.read_add_innervmstubin(VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2_read_add),
.innervmstubin(VMS_F1D5PHI2X2n2_TE_F1D5PHI2X2_F2D5PHI2X2),
.stubpairout(TE_F1D5PHI2X2_F2D5PHI2X2_SP_F1D5PHI2X2_F2D5PHI2X2),
.valid_data(TE_F1D5PHI2X2_F2D5PHI2X2_SP_F1D5PHI2X2_F2D5PHI2X2_wr_en),
.start(VMS_F2D5PHI2X2n3_start),
.done(TE_F1D5PHI2X2_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI3X2_F2D5PHI2X2_phi.txt","TETable_TE_F1D5PHI3X2_F2D5PHI2X2_z.txt",1'b0) TE_F1D5PHI3X2_F2D5PHI2X2(
.number_in_outervmstubin(VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2_number),
.read_add_outervmstubin(VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2_read_add),
.outervmstubin(VMS_F2D5PHI2X2n4_TE_F1D5PHI3X2_F2D5PHI2X2),
.number_in_innervmstubin(VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2_number),
.read_add_innervmstubin(VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2_read_add),
.innervmstubin(VMS_F1D5PHI3X2n1_TE_F1D5PHI3X2_F2D5PHI2X2),
.stubpairout(TE_F1D5PHI3X2_F2D5PHI2X2_SP_F1D5PHI3X2_F2D5PHI2X2),
.valid_data(TE_F1D5PHI3X2_F2D5PHI2X2_SP_F1D5PHI3X2_F2D5PHI2X2_wr_en),
.start(VMS_F2D5PHI2X2n4_start),
.done(TE_F1D5PHI3X2_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI3X2_F2D5PHI3X2_phi.txt","TETable_TE_F1D5PHI3X2_F2D5PHI3X2_z.txt",1'b0) TE_F1D5PHI3X2_F2D5PHI3X2(
.number_in_outervmstubin(VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2_number),
.read_add_outervmstubin(VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2_read_add),
.outervmstubin(VMS_F2D5PHI3X2n3_TE_F1D5PHI3X2_F2D5PHI3X2),
.number_in_innervmstubin(VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2_number),
.read_add_innervmstubin(VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2_read_add),
.innervmstubin(VMS_F1D5PHI3X2n2_TE_F1D5PHI3X2_F2D5PHI3X2),
.stubpairout(TE_F1D5PHI3X2_F2D5PHI3X2_SP_F1D5PHI3X2_F2D5PHI3X2),
.valid_data(TE_F1D5PHI3X2_F2D5PHI3X2_SP_F1D5PHI3X2_F2D5PHI3X2_wr_en),
.start(VMS_F2D5PHI3X2n3_start),
.done(TE_F1D5PHI3X2_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F1D5PHI4X2_F2D5PHI3X2_phi.txt","TETable_TE_F1D5PHI4X2_F2D5PHI3X2_z.txt",1'b0) TE_F1D5PHI4X2_F2D5PHI3X2(
.number_in_outervmstubin(VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2_number),
.read_add_outervmstubin(VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2_read_add),
.outervmstubin(VMS_F2D5PHI3X2n4_TE_F1D5PHI4X2_F2D5PHI3X2),
.number_in_innervmstubin(VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2_number),
.read_add_innervmstubin(VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2_read_add),
.innervmstubin(VMS_F1D5PHI4X2n1_TE_F1D5PHI4X2_F2D5PHI3X2),
.stubpairout(TE_F1D5PHI4X2_F2D5PHI3X2_SP_F1D5PHI4X2_F2D5PHI3X2),
.valid_data(TE_F1D5PHI4X2_F2D5PHI3X2_SP_F1D5PHI4X2_F2D5PHI3X2_wr_en),
.start(VMS_F2D5PHI3X2n4_start),
.done(TE_F1D5PHI4X2_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI1X1_F4D5PHI1X1_phi.txt","TETable_TE_F3D5PHI1X1_F4D5PHI1X1_z.txt",1'b0) TE_F3D5PHI1X1_F4D5PHI1X1(
.number_in_innervmstubin(VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_number),
.read_add_innervmstubin(VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_read_add),
.innervmstubin(VMS_F3D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1),
.number_in_outervmstubin(VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_number),
.read_add_outervmstubin(VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1_read_add),
.outervmstubin(VMS_F4D5PHI1X1n1_TE_F3D5PHI1X1_F4D5PHI1X1),
.stubpairout(TE_F3D5PHI1X1_F4D5PHI1X1_SP_F3D5PHI1X1_F4D5PHI1X1),
.valid_data(TE_F3D5PHI1X1_F4D5PHI1X1_SP_F3D5PHI1X1_F4D5PHI1X1_wr_en),
.start(VMS_F3D5PHI1X1n1_start),
.done(TE_F3D5PHI1X1_F4D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI2X1_F4D5PHI1X1_phi.txt","TETable_TE_F3D5PHI2X1_F4D5PHI1X1_z.txt",1'b0) TE_F3D5PHI2X1_F4D5PHI1X1(
.number_in_outervmstubin(VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1_number),
.read_add_outervmstubin(VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1_read_add),
.outervmstubin(VMS_F4D5PHI1X1n2_TE_F3D5PHI2X1_F4D5PHI1X1),
.number_in_innervmstubin(VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1_number),
.read_add_innervmstubin(VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1_read_add),
.innervmstubin(VMS_F3D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI1X1),
.stubpairout(TE_F3D5PHI2X1_F4D5PHI1X1_SP_F3D5PHI2X1_F4D5PHI1X1),
.valid_data(TE_F3D5PHI2X1_F4D5PHI1X1_SP_F3D5PHI2X1_F4D5PHI1X1_wr_en),
.start(VMS_F4D5PHI1X1n2_start),
.done(TE_F3D5PHI2X1_F4D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI2X1_F4D5PHI2X1_phi.txt","TETable_TE_F3D5PHI2X1_F4D5PHI2X1_z.txt",1'b0) TE_F3D5PHI2X1_F4D5PHI2X1(
.number_in_innervmstubin(VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1_number),
.read_add_innervmstubin(VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1_read_add),
.innervmstubin(VMS_F3D5PHI2X1n2_TE_F3D5PHI2X1_F4D5PHI2X1),
.number_in_outervmstubin(VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1_number),
.read_add_outervmstubin(VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1_read_add),
.outervmstubin(VMS_F4D5PHI2X1n1_TE_F3D5PHI2X1_F4D5PHI2X1),
.stubpairout(TE_F3D5PHI2X1_F4D5PHI2X1_SP_F3D5PHI2X1_F4D5PHI2X1),
.valid_data(TE_F3D5PHI2X1_F4D5PHI2X1_SP_F3D5PHI2X1_F4D5PHI2X1_wr_en),
.start(VMS_F3D5PHI2X1n2_start),
.done(TE_F3D5PHI2X1_F4D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI3X1_F4D5PHI2X1_phi.txt","TETable_TE_F3D5PHI3X1_F4D5PHI2X1_z.txt",1'b0) TE_F3D5PHI3X1_F4D5PHI2X1(
.number_in_outervmstubin(VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1_number),
.read_add_outervmstubin(VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1_read_add),
.outervmstubin(VMS_F4D5PHI2X1n2_TE_F3D5PHI3X1_F4D5PHI2X1),
.number_in_innervmstubin(VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1_number),
.read_add_innervmstubin(VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1_read_add),
.innervmstubin(VMS_F3D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI2X1),
.stubpairout(TE_F3D5PHI3X1_F4D5PHI2X1_SP_F3D5PHI3X1_F4D5PHI2X1),
.valid_data(TE_F3D5PHI3X1_F4D5PHI2X1_SP_F3D5PHI3X1_F4D5PHI2X1_wr_en),
.start(VMS_F4D5PHI2X1n2_start),
.done(TE_F3D5PHI3X1_F4D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI3X1_F4D5PHI3X1_phi.txt","TETable_TE_F3D5PHI3X1_F4D5PHI3X1_z.txt",1'b0) TE_F3D5PHI3X1_F4D5PHI3X1(
.number_in_innervmstubin(VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1_number),
.read_add_innervmstubin(VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1_read_add),
.innervmstubin(VMS_F3D5PHI3X1n2_TE_F3D5PHI3X1_F4D5PHI3X1),
.number_in_outervmstubin(VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1_number),
.read_add_outervmstubin(VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1_read_add),
.outervmstubin(VMS_F4D5PHI3X1n1_TE_F3D5PHI3X1_F4D5PHI3X1),
.stubpairout(TE_F3D5PHI3X1_F4D5PHI3X1_SP_F3D5PHI3X1_F4D5PHI3X1),
.valid_data(TE_F3D5PHI3X1_F4D5PHI3X1_SP_F3D5PHI3X1_F4D5PHI3X1_wr_en),
.start(VMS_F3D5PHI3X1n2_start),
.done(TE_F3D5PHI3X1_F4D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI4X1_F4D5PHI3X1_phi.txt","TETable_TE_F3D5PHI4X1_F4D5PHI3X1_z.txt",1'b0) TE_F3D5PHI4X1_F4D5PHI3X1(
.number_in_outervmstubin(VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1_number),
.read_add_outervmstubin(VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1_read_add),
.outervmstubin(VMS_F4D5PHI3X1n2_TE_F3D5PHI4X1_F4D5PHI3X1),
.number_in_innervmstubin(VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1_number),
.read_add_innervmstubin(VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1_read_add),
.innervmstubin(VMS_F3D5PHI4X1n1_TE_F3D5PHI4X1_F4D5PHI3X1),
.stubpairout(TE_F3D5PHI4X1_F4D5PHI3X1_SP_F3D5PHI4X1_F4D5PHI3X1),
.valid_data(TE_F3D5PHI4X1_F4D5PHI3X1_SP_F3D5PHI4X1_F4D5PHI3X1_wr_en),
.start(VMS_F4D5PHI3X1n2_start),
.done(TE_F3D5PHI4X1_F4D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI1X1_F4D5PHI1X2_phi.txt","TETable_TE_F3D5PHI1X1_F4D5PHI1X2_z.txt",1'b0) TE_F3D5PHI1X1_F4D5PHI1X2(
.number_in_innervmstubin(VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2_number),
.read_add_innervmstubin(VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2_read_add),
.innervmstubin(VMS_F3D5PHI1X1n2_TE_F3D5PHI1X1_F4D5PHI1X2),
.number_in_outervmstubin(VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2_number),
.read_add_outervmstubin(VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2_read_add),
.outervmstubin(VMS_F4D5PHI1X2n1_TE_F3D5PHI1X1_F4D5PHI1X2),
.stubpairout(TE_F3D5PHI1X1_F4D5PHI1X2_SP_F3D5PHI1X1_F4D5PHI1X2),
.valid_data(TE_F3D5PHI1X1_F4D5PHI1X2_SP_F3D5PHI1X1_F4D5PHI1X2_wr_en),
.start(VMS_F3D5PHI1X1n2_start),
.done(TE_F3D5PHI1X1_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI2X1_F4D5PHI1X2_phi.txt","TETable_TE_F3D5PHI2X1_F4D5PHI1X2_z.txt",1'b0) TE_F3D5PHI2X1_F4D5PHI1X2(
.number_in_innervmstubin(VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2_number),
.read_add_innervmstubin(VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2_read_add),
.innervmstubin(VMS_F3D5PHI2X1n3_TE_F3D5PHI2X1_F4D5PHI1X2),
.number_in_outervmstubin(VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2_number),
.read_add_outervmstubin(VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2_read_add),
.outervmstubin(VMS_F4D5PHI1X2n2_TE_F3D5PHI2X1_F4D5PHI1X2),
.stubpairout(TE_F3D5PHI2X1_F4D5PHI1X2_SP_F3D5PHI2X1_F4D5PHI1X2),
.valid_data(TE_F3D5PHI2X1_F4D5PHI1X2_SP_F3D5PHI2X1_F4D5PHI1X2_wr_en),
.start(VMS_F3D5PHI2X1n3_start),
.done(TE_F3D5PHI2X1_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI2X1_F4D5PHI2X2_phi.txt","TETable_TE_F3D5PHI2X1_F4D5PHI2X2_z.txt",1'b0) TE_F3D5PHI2X1_F4D5PHI2X2(
.number_in_innervmstubin(VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2_number),
.read_add_innervmstubin(VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2_read_add),
.innervmstubin(VMS_F3D5PHI2X1n4_TE_F3D5PHI2X1_F4D5PHI2X2),
.number_in_outervmstubin(VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2_number),
.read_add_outervmstubin(VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2_read_add),
.outervmstubin(VMS_F4D5PHI2X2n1_TE_F3D5PHI2X1_F4D5PHI2X2),
.stubpairout(TE_F3D5PHI2X1_F4D5PHI2X2_SP_F3D5PHI2X1_F4D5PHI2X2),
.valid_data(TE_F3D5PHI2X1_F4D5PHI2X2_SP_F3D5PHI2X1_F4D5PHI2X2_wr_en),
.start(VMS_F3D5PHI2X1n4_start),
.done(TE_F3D5PHI2X1_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI3X1_F4D5PHI2X2_phi.txt","TETable_TE_F3D5PHI3X1_F4D5PHI2X2_z.txt",1'b0) TE_F3D5PHI3X1_F4D5PHI2X2(
.number_in_innervmstubin(VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2_number),
.read_add_innervmstubin(VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2_read_add),
.innervmstubin(VMS_F3D5PHI3X1n3_TE_F3D5PHI3X1_F4D5PHI2X2),
.number_in_outervmstubin(VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2_number),
.read_add_outervmstubin(VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2_read_add),
.outervmstubin(VMS_F4D5PHI2X2n2_TE_F3D5PHI3X1_F4D5PHI2X2),
.stubpairout(TE_F3D5PHI3X1_F4D5PHI2X2_SP_F3D5PHI3X1_F4D5PHI2X2),
.valid_data(TE_F3D5PHI3X1_F4D5PHI2X2_SP_F3D5PHI3X1_F4D5PHI2X2_wr_en),
.start(VMS_F3D5PHI3X1n3_start),
.done(TE_F3D5PHI3X1_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI3X1_F4D5PHI3X2_phi.txt","TETable_TE_F3D5PHI3X1_F4D5PHI3X2_z.txt",1'b0) TE_F3D5PHI3X1_F4D5PHI3X2(
.number_in_innervmstubin(VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2_number),
.read_add_innervmstubin(VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2_read_add),
.innervmstubin(VMS_F3D5PHI3X1n4_TE_F3D5PHI3X1_F4D5PHI3X2),
.number_in_outervmstubin(VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2_number),
.read_add_outervmstubin(VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2_read_add),
.outervmstubin(VMS_F4D5PHI3X2n1_TE_F3D5PHI3X1_F4D5PHI3X2),
.stubpairout(TE_F3D5PHI3X1_F4D5PHI3X2_SP_F3D5PHI3X1_F4D5PHI3X2),
.valid_data(TE_F3D5PHI3X1_F4D5PHI3X2_SP_F3D5PHI3X1_F4D5PHI3X2_wr_en),
.start(VMS_F3D5PHI3X1n4_start),
.done(TE_F3D5PHI3X1_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI4X1_F4D5PHI3X2_phi.txt","TETable_TE_F3D5PHI4X1_F4D5PHI3X2_z.txt",1'b0) TE_F3D5PHI4X1_F4D5PHI3X2(
.number_in_innervmstubin(VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2_number),
.read_add_innervmstubin(VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2_read_add),
.innervmstubin(VMS_F3D5PHI4X1n2_TE_F3D5PHI4X1_F4D5PHI3X2),
.number_in_outervmstubin(VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2_number),
.read_add_outervmstubin(VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2_read_add),
.outervmstubin(VMS_F4D5PHI3X2n2_TE_F3D5PHI4X1_F4D5PHI3X2),
.stubpairout(TE_F3D5PHI4X1_F4D5PHI3X2_SP_F3D5PHI4X1_F4D5PHI3X2),
.valid_data(TE_F3D5PHI4X1_F4D5PHI3X2_SP_F3D5PHI4X1_F4D5PHI3X2_wr_en),
.start(VMS_F3D5PHI4X1n2_start),
.done(TE_F3D5PHI4X1_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI1X2_F4D5PHI1X2_phi.txt","TETable_TE_F3D5PHI1X2_F4D5PHI1X2_z.txt",1'b0) TE_F3D5PHI1X2_F4D5PHI1X2(
.number_in_outervmstubin(VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2_number),
.read_add_outervmstubin(VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2_read_add),
.outervmstubin(VMS_F4D5PHI1X2n3_TE_F3D5PHI1X2_F4D5PHI1X2),
.number_in_innervmstubin(VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2_number),
.read_add_innervmstubin(VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2_read_add),
.innervmstubin(VMS_F3D5PHI1X2n1_TE_F3D5PHI1X2_F4D5PHI1X2),
.stubpairout(TE_F3D5PHI1X2_F4D5PHI1X2_SP_F3D5PHI1X2_F4D5PHI1X2),
.valid_data(TE_F3D5PHI1X2_F4D5PHI1X2_SP_F3D5PHI1X2_F4D5PHI1X2_wr_en),
.start(VMS_F4D5PHI1X2n3_start),
.done(TE_F3D5PHI1X2_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI2X2_F4D5PHI1X2_phi.txt","TETable_TE_F3D5PHI2X2_F4D5PHI1X2_z.txt",1'b0) TE_F3D5PHI2X2_F4D5PHI1X2(
.number_in_outervmstubin(VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2_number),
.read_add_outervmstubin(VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2_read_add),
.outervmstubin(VMS_F4D5PHI1X2n4_TE_F3D5PHI2X2_F4D5PHI1X2),
.number_in_innervmstubin(VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2_number),
.read_add_innervmstubin(VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2_read_add),
.innervmstubin(VMS_F3D5PHI2X2n1_TE_F3D5PHI2X2_F4D5PHI1X2),
.stubpairout(TE_F3D5PHI2X2_F4D5PHI1X2_SP_F3D5PHI2X2_F4D5PHI1X2),
.valid_data(TE_F3D5PHI2X2_F4D5PHI1X2_SP_F3D5PHI2X2_F4D5PHI1X2_wr_en),
.start(VMS_F4D5PHI1X2n4_start),
.done(TE_F3D5PHI2X2_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI2X2_F4D5PHI2X2_phi.txt","TETable_TE_F3D5PHI2X2_F4D5PHI2X2_z.txt",1'b0) TE_F3D5PHI2X2_F4D5PHI2X2(
.number_in_outervmstubin(VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2_number),
.read_add_outervmstubin(VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2_read_add),
.outervmstubin(VMS_F4D5PHI2X2n3_TE_F3D5PHI2X2_F4D5PHI2X2),
.number_in_innervmstubin(VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2_number),
.read_add_innervmstubin(VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2_read_add),
.innervmstubin(VMS_F3D5PHI2X2n2_TE_F3D5PHI2X2_F4D5PHI2X2),
.stubpairout(TE_F3D5PHI2X2_F4D5PHI2X2_SP_F3D5PHI2X2_F4D5PHI2X2),
.valid_data(TE_F3D5PHI2X2_F4D5PHI2X2_SP_F3D5PHI2X2_F4D5PHI2X2_wr_en),
.start(VMS_F4D5PHI2X2n3_start),
.done(TE_F3D5PHI2X2_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI3X2_F4D5PHI2X2_phi.txt","TETable_TE_F3D5PHI3X2_F4D5PHI2X2_z.txt",1'b0) TE_F3D5PHI3X2_F4D5PHI2X2(
.number_in_outervmstubin(VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2_number),
.read_add_outervmstubin(VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2_read_add),
.outervmstubin(VMS_F4D5PHI2X2n4_TE_F3D5PHI3X2_F4D5PHI2X2),
.number_in_innervmstubin(VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2_number),
.read_add_innervmstubin(VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2_read_add),
.innervmstubin(VMS_F3D5PHI3X2n1_TE_F3D5PHI3X2_F4D5PHI2X2),
.stubpairout(TE_F3D5PHI3X2_F4D5PHI2X2_SP_F3D5PHI3X2_F4D5PHI2X2),
.valid_data(TE_F3D5PHI3X2_F4D5PHI2X2_SP_F3D5PHI3X2_F4D5PHI2X2_wr_en),
.start(VMS_F4D5PHI2X2n4_start),
.done(TE_F3D5PHI3X2_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI3X2_F4D5PHI3X2_phi.txt","TETable_TE_F3D5PHI3X2_F4D5PHI3X2_z.txt",1'b0) TE_F3D5PHI3X2_F4D5PHI3X2(
.number_in_outervmstubin(VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2_number),
.read_add_outervmstubin(VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2_read_add),
.outervmstubin(VMS_F4D5PHI3X2n3_TE_F3D5PHI3X2_F4D5PHI3X2),
.number_in_innervmstubin(VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2_number),
.read_add_innervmstubin(VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2_read_add),
.innervmstubin(VMS_F3D5PHI3X2n2_TE_F3D5PHI3X2_F4D5PHI3X2),
.stubpairout(TE_F3D5PHI3X2_F4D5PHI3X2_SP_F3D5PHI3X2_F4D5PHI3X2),
.valid_data(TE_F3D5PHI3X2_F4D5PHI3X2_SP_F3D5PHI3X2_F4D5PHI3X2_wr_en),
.start(VMS_F4D5PHI3X2n3_start),
.done(TE_F3D5PHI3X2_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_F3D5PHI4X2_F4D5PHI3X2_phi.txt","TETable_TE_F3D5PHI4X2_F4D5PHI3X2_z.txt",1'b0) TE_F3D5PHI4X2_F4D5PHI3X2(
.number_in_outervmstubin(VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2_number),
.read_add_outervmstubin(VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2_read_add),
.outervmstubin(VMS_F4D5PHI3X2n4_TE_F3D5PHI4X2_F4D5PHI3X2),
.number_in_innervmstubin(VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2_number),
.read_add_innervmstubin(VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2_read_add),
.innervmstubin(VMS_F3D5PHI4X2n1_TE_F3D5PHI4X2_F4D5PHI3X2),
.stubpairout(TE_F3D5PHI4X2_F4D5PHI3X2_SP_F3D5PHI4X2_F4D5PHI3X2),
.valid_data(TE_F3D5PHI4X2_F4D5PHI3X2_SP_F3D5PHI4X2_F4D5PHI3X2_wr_en),
.start(VMS_F4D5PHI3X2n4_start),
.done(TE_F3D5PHI4X2_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(0),.InvR_FILE("InvRTable_TC_F1D5F2D5.dat"),.InvT_FILE("InvTTable_TC_F1D5F2D5.dat"),.TC_index(4'b0100)) TC_F1D5F2D5(
.number_in_stubpair1in(SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5_number),
.read_add_stubpair1in(SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5_read_add),
.stubpair1in(SP_F1D5PHI1X1_F2D5PHI1X1_TC_F1D5F2D5),
.number_in_stubpair2in(SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5_number),
.read_add_stubpair2in(SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5_read_add),
.stubpair2in(SP_F1D5PHI2X1_F2D5PHI1X1_TC_F1D5F2D5),
.number_in_stubpair3in(SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5_number),
.read_add_stubpair3in(SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5_read_add),
.stubpair3in(SP_F1D5PHI2X1_F2D5PHI2X1_TC_F1D5F2D5),
.number_in_stubpair4in(SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5_number),
.read_add_stubpair4in(SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5_read_add),
.stubpair4in(SP_F1D5PHI3X1_F2D5PHI2X1_TC_F1D5F2D5),
.number_in_stubpair5in(SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5_number),
.read_add_stubpair5in(SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5_read_add),
.stubpair5in(SP_F1D5PHI3X1_F2D5PHI3X1_TC_F1D5F2D5),
.number_in_stubpair6in(SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5_number),
.read_add_stubpair6in(SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5_read_add),
.stubpair6in(SP_F1D5PHI4X1_F2D5PHI3X1_TC_F1D5F2D5),
.number_in_stubpair7in(SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5_number),
.read_add_stubpair7in(SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5_read_add),
.stubpair7in(SP_F1D5PHI1X1_F2D5PHI1X2_TC_F1D5F2D5),
.number_in_stubpair8in(SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5_number),
.read_add_stubpair8in(SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5_read_add),
.stubpair8in(SP_F1D5PHI2X1_F2D5PHI1X2_TC_F1D5F2D5),
.number_in_stubpair9in(SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5_number),
.read_add_stubpair9in(SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5_read_add),
.stubpair9in(SP_F1D5PHI2X1_F2D5PHI2X2_TC_F1D5F2D5),
.number_in_stubpair10in(SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5_number),
.read_add_stubpair10in(SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5_read_add),
.stubpair10in(SP_F1D5PHI3X1_F2D5PHI2X2_TC_F1D5F2D5),
.number_in_stubpair11in(SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5_number),
.read_add_stubpair11in(SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5_read_add),
.stubpair11in(SP_F1D5PHI3X1_F2D5PHI3X2_TC_F1D5F2D5),
.number_in_stubpair12in(SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5_number),
.read_add_stubpair12in(SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5_read_add),
.stubpair12in(SP_F1D5PHI4X1_F2D5PHI3X2_TC_F1D5F2D5),
.number_in_stubpair13in(SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5_number),
.read_add_stubpair13in(SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5_read_add),
.stubpair13in(SP_F1D5PHI1X2_F2D5PHI1X2_TC_F1D5F2D5),
.number_in_stubpair14in(SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5_number),
.read_add_stubpair14in(SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5_read_add),
.stubpair14in(SP_F1D5PHI2X2_F2D5PHI1X2_TC_F1D5F2D5),
.number_in_stubpair15in(SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5_number),
.read_add_stubpair15in(SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5_read_add),
.stubpair15in(SP_F1D5PHI2X2_F2D5PHI2X2_TC_F1D5F2D5),
.number_in_stubpair16in(SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5_number),
.read_add_stubpair16in(SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5_read_add),
.stubpair16in(SP_F1D5PHI3X2_F2D5PHI2X2_TC_F1D5F2D5),
.number_in_stubpair17in(SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5_number),
.read_add_stubpair17in(SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5_read_add),
.stubpair17in(SP_F1D5PHI3X2_F2D5PHI3X2_TC_F1D5F2D5),
.number_in_stubpair18in(SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5_number),
.read_add_stubpair18in(SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5_read_add),
.stubpair18in(SP_F1D5PHI4X2_F2D5PHI3X2_TC_F1D5F2D5),
.read_add_outerallstubin(AS_F2D5n1_TC_F1D5F2D5_read_add),
.outerallstubin(AS_F2D5n1_TC_F1D5F2D5),
.read_add_innerallstubin(AS_F1D5n1_TC_F1D5F2D5_read_add),
.innerallstubin(AS_F1D5n1_TC_F1D5F2D5),
.projoutToPlus_F5(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F5),
.projoutToPlus_F3(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F3),
.projoutToPlus_F4(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F4),
.projoutToMinus_F5(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F5),
.projoutToMinus_F3(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F3),
.projoutToMinus_F4(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F4),
.projout_F3D5(TC_F1D5F2D5_TPROJ_F1D5F2D5_F3D5),
.projout_F4D5(TC_F1D5F2D5_TPROJ_F1D5F2D5_F4D5),
.projout_F5D5(TC_F1D5F2D5_TPROJ_F1D5F2D5_F5D5),
.trackpar(TC_F1D5F2D5_TPAR_F1D5F2D5),
.valid_projoutToPlus_F5(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F5_wr_en),
.valid_projoutToPlus_F3(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F3_wr_en),
.valid_projoutToPlus_F4(TC_F1D5F2D5_TPROJ_ToPlus_F1D5F2D5_F4_wr_en),
.valid_projoutToMinus_F5(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F5_wr_en),
.valid_projoutToMinus_F3(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F3_wr_en),
.valid_projoutToMinus_F4(TC_F1D5F2D5_TPROJ_ToMinus_F1D5F2D5_F4_wr_en),
.valid_projout_F3D5(TC_F1D5F2D5_TPROJ_F1D5F2D5_F3D5_wr_en),
.valid_projout_F4D5(TC_F1D5F2D5_TPROJ_F1D5F2D5_F4D5_wr_en),
.valid_projout_F5D5(TC_F1D5F2D5_TPROJ_F1D5F2D5_F5D5_wr_en),
.valid_trackpar(TC_F1D5F2D5_TPAR_F1D5F2D5_wr_en),
.done_proj(TC_F1D5F2D5_proj_start),
.start(SP_F1D5PHI1X1_F2D5PHI1X1_start),
.done(TC_F1D5F2D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(0),.InvR_FILE("InvRTable_TC_F3D5F4D5.dat"),.InvT_FILE("InvTTable_TC_F3D5F4D5.dat"),.TC_index(4'b0100)) TC_F3D5F4D5(
.number_in_stubpair1in(SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5_number),
.read_add_stubpair1in(SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5_read_add),
.stubpair1in(SP_F3D5PHI1X1_F4D5PHI1X1_TC_F3D5F4D5),
.number_in_stubpair2in(SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5_number),
.read_add_stubpair2in(SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5_read_add),
.stubpair2in(SP_F3D5PHI2X1_F4D5PHI1X1_TC_F3D5F4D5),
.number_in_stubpair3in(SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5_number),
.read_add_stubpair3in(SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5_read_add),
.stubpair3in(SP_F3D5PHI2X1_F4D5PHI2X1_TC_F3D5F4D5),
.number_in_stubpair4in(SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5_number),
.read_add_stubpair4in(SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5_read_add),
.stubpair4in(SP_F3D5PHI3X1_F4D5PHI2X1_TC_F3D5F4D5),
.number_in_stubpair5in(SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5_number),
.read_add_stubpair5in(SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5_read_add),
.stubpair5in(SP_F3D5PHI3X1_F4D5PHI3X1_TC_F3D5F4D5),
.number_in_stubpair6in(SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5_number),
.read_add_stubpair6in(SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5_read_add),
.stubpair6in(SP_F3D5PHI4X1_F4D5PHI3X1_TC_F3D5F4D5),
.number_in_stubpair7in(SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5_number),
.read_add_stubpair7in(SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5_read_add),
.stubpair7in(SP_F3D5PHI1X1_F4D5PHI1X2_TC_F3D5F4D5),
.number_in_stubpair8in(SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5_number),
.read_add_stubpair8in(SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5_read_add),
.stubpair8in(SP_F3D5PHI2X1_F4D5PHI1X2_TC_F3D5F4D5),
.number_in_stubpair9in(SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5_number),
.read_add_stubpair9in(SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5_read_add),
.stubpair9in(SP_F3D5PHI2X1_F4D5PHI2X2_TC_F3D5F4D5),
.number_in_stubpair10in(SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5_number),
.read_add_stubpair10in(SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5_read_add),
.stubpair10in(SP_F3D5PHI3X1_F4D5PHI2X2_TC_F3D5F4D5),
.number_in_stubpair11in(SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5_number),
.read_add_stubpair11in(SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5_read_add),
.stubpair11in(SP_F3D5PHI3X1_F4D5PHI3X2_TC_F3D5F4D5),
.number_in_stubpair12in(SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5_number),
.read_add_stubpair12in(SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5_read_add),
.stubpair12in(SP_F3D5PHI4X1_F4D5PHI3X2_TC_F3D5F4D5),
.number_in_stubpair13in(SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5_number),
.read_add_stubpair13in(SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5_read_add),
.stubpair13in(SP_F3D5PHI1X2_F4D5PHI1X2_TC_F3D5F4D5),
.number_in_stubpair14in(SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5_number),
.read_add_stubpair14in(SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5_read_add),
.stubpair14in(SP_F3D5PHI2X2_F4D5PHI1X2_TC_F3D5F4D5),
.number_in_stubpair15in(SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5_number),
.read_add_stubpair15in(SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5_read_add),
.stubpair15in(SP_F3D5PHI2X2_F4D5PHI2X2_TC_F3D5F4D5),
.number_in_stubpair16in(SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5_number),
.read_add_stubpair16in(SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5_read_add),
.stubpair16in(SP_F3D5PHI3X2_F4D5PHI2X2_TC_F3D5F4D5),
.number_in_stubpair17in(SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5_number),
.read_add_stubpair17in(SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5_read_add),
.stubpair17in(SP_F3D5PHI3X2_F4D5PHI3X2_TC_F3D5F4D5),
.number_in_stubpair18in(SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5_number),
.read_add_stubpair18in(SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5_read_add),
.stubpair18in(SP_F3D5PHI4X2_F4D5PHI3X2_TC_F3D5F4D5),
.read_add_outerallstubin(AS_F4D5n1_TC_F3D5F4D5_read_add),
.outerallstubin(AS_F4D5n1_TC_F3D5F4D5),
.read_add_innerallstubin(AS_F3D5n1_TC_F3D5F4D5_read_add),
.innerallstubin(AS_F3D5n1_TC_F3D5F4D5),
.projoutToPlus_F5(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F5),
.projoutToPlus_F2(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F2),
.projoutToPlus_F1(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F1),
.projoutToMinus_F5(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F5),
.projoutToMinus_F2(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F2),
.projoutToMinus_F1(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F1),
.projout_F1D5(TC_F3D5F4D5_TPROJ_F3D5F4D5_F1D5),
.projout_F2D5(TC_F3D5F4D5_TPROJ_F3D5F4D5_F2D5),
.projout_F5D5(TC_F3D5F4D5_TPROJ_F3D5F4D5_F5D5),
.trackpar(TC_F3D5F4D5_TPAR_F3D5F4D5),
.valid_projoutToPlus_F5(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F5_wr_en),
.valid_projoutToPlus_F2(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F2_wr_en),
.valid_projoutToPlus_F1(TC_F3D5F4D5_TPROJ_ToPlus_F3D5F4D5_F1_wr_en),
.valid_projoutToMinus_F5(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F5_wr_en),
.valid_projoutToMinus_F2(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F2_wr_en),
.valid_projoutToMinus_F1(TC_F3D5F4D5_TPROJ_ToMinus_F3D5F4D5_F1_wr_en),
.valid_projout_F1D5(TC_F3D5F4D5_TPROJ_F3D5F4D5_F1D5_wr_en),
.valid_projout_F2D5(TC_F3D5F4D5_TPROJ_F3D5F4D5_F2D5_wr_en),
.valid_projout_F5D5(TC_F3D5F4D5_TPROJ_F3D5F4D5_F5D5_wr_en),
.valid_trackpar(TC_F3D5F4D5_TPAR_F3D5F4D5_wr_en),
.done_proj(TC_F3D5F4D5_proj_start),
.start(SP_F3D5PHI1X1_F4D5PHI1X1_start),
.done(TC_F3D5F4D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b0,1'b0) PRD_F3D5_F1F2(
.number_in_proj1in(TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2_number),
.read_add_proj1in(TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2_read_add),
.proj1in(TPROJ_FromPlus_F3D5_F1F2_PRD_F3D5_F1F2),
.number_in_proj2in(TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2_number),
.read_add_proj2in(TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2_read_add),
.proj2in(TPROJ_FromMinus_F3D5_F1F2_PRD_F3D5_F1F2),
.number_in_proj3in(TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2_number),
.read_add_proj3in(TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2_read_add),
.proj3in(TPROJ_F1D5F2D5_F3D5_PRD_F3D5_F1F2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X1),
.vmprojoutPHI1X2(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X2),
.vmprojoutPHI2X1(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X1),
.vmprojoutPHI2X2(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X2),
.vmprojoutPHI3X1(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X1),
.vmprojoutPHI3X2(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X2),
.vmprojoutPHI4X1(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X1),
.vmprojoutPHI4X2(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X2),
.allprojout(PRD_F3D5_F1F2_AP_F1F2_F3D5),
.valid_data(PRD_F3D5_F1F2_AP_F1F2_F3D5_wr_en),
.vmprojoutPHI1X1_wr_en(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PRD_F3D5_F1F2_VMPROJ_F1F2_F3D5PHI4X2_wr_en),
.start(TPROJ_FromPlus_F3D5_F1F2_start),
.done(PRD_F3D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0,1'b0) PRD_F4D5_F1F2(
.number_in_proj1in(TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2_number),
.read_add_proj1in(TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2_read_add),
.proj1in(TPROJ_FromPlus_F4D5_F1F2_PRD_F4D5_F1F2),
.number_in_proj2in(TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2_number),
.read_add_proj2in(TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2_read_add),
.proj2in(TPROJ_FromMinus_F4D5_F1F2_PRD_F4D5_F1F2),
.number_in_proj3in(TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2_number),
.read_add_proj3in(TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2_read_add),
.proj3in(TPROJ_F1D5F2D5_F4D5_PRD_F4D5_F1F2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X1),
.vmprojoutPHI1X2(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X2),
.vmprojoutPHI2X1(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X1),
.vmprojoutPHI2X2(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X2),
.vmprojoutPHI3X1(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X1),
.vmprojoutPHI3X2(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X2),
.allprojout(PRD_F4D5_F1F2_AP_F1F2_F4D5),
.valid_data(PRD_F4D5_F1F2_AP_F1F2_F4D5_wr_en),
.vmprojoutPHI1X1_wr_en(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PRD_F4D5_F1F2_VMPROJ_F1F2_F4D5PHI3X2_wr_en),
.start(TPROJ_FromPlus_F4D5_F1F2_start),
.done(PRD_F4D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b0,1'b0) PRD_F5D5_F1F2(
.number_in_proj1in(TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2_number),
.read_add_proj1in(TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2_read_add),
.proj1in(TPROJ_FromPlus_F5D5_F1F2_PRD_F5D5_F1F2),
.number_in_proj2in(TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2_number),
.read_add_proj2in(TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2_read_add),
.proj2in(TPROJ_FromMinus_F5D5_F1F2_PRD_F5D5_F1F2),
.number_in_proj3in(TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2_number),
.read_add_proj3in(TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2_read_add),
.proj3in(TPROJ_F1D5F2D5_F5D5_PRD_F5D5_F1F2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X1),
.vmprojoutPHI1X2(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X2),
.vmprojoutPHI2X1(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X1),
.vmprojoutPHI2X2(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X2),
.vmprojoutPHI3X1(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X1),
.vmprojoutPHI3X2(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X2),
.vmprojoutPHI4X1(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X1),
.vmprojoutPHI4X2(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X2),
.allprojout(PRD_F5D5_F1F2_AP_F1F2_F5D5),
.valid_data(PRD_F5D5_F1F2_AP_F1F2_F5D5_wr_en),
.vmprojoutPHI1X1_wr_en(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PRD_F5D5_F1F2_VMPROJ_F1F2_F5D5PHI4X2_wr_en),
.start(TPROJ_FromPlus_F5D5_F1F2_start),
.done(PRD_F5D5_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b0,1'b0) PRD_F1D5_F3F4(
.number_in_proj1in(TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4_number),
.read_add_proj1in(TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4_read_add),
.proj1in(TPROJ_FromPlus_F1D5_F3F4_PRD_F1D5_F3F4),
.number_in_proj2in(TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4_number),
.read_add_proj2in(TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4_read_add),
.proj2in(TPROJ_FromMinus_F1D5_F3F4_PRD_F1D5_F3F4),
.number_in_proj3in(TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4_number),
.read_add_proj3in(TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4_read_add),
.proj3in(TPROJ_F3D5F4D5_F1D5_PRD_F1D5_F3F4),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X1),
.vmprojoutPHI1X2(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X2),
.vmprojoutPHI2X1(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X1),
.vmprojoutPHI2X2(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X2),
.vmprojoutPHI3X1(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X1),
.vmprojoutPHI3X2(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X2),
.vmprojoutPHI4X1(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X1),
.vmprojoutPHI4X2(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X2),
.allprojout(PRD_F1D5_F3F4_AP_F3F4_F1D5),
.valid_data(PRD_F1D5_F3F4_AP_F3F4_F1D5_wr_en),
.vmprojoutPHI1X1_wr_en(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PRD_F1D5_F3F4_VMPROJ_F3F4_F1D5PHI4X2_wr_en),
.start(TPROJ_FromPlus_F1D5_F3F4_start),
.done(PRD_F1D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0,1'b0) PRD_F2D5_F3F4(
.number_in_proj1in(TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4_number),
.read_add_proj1in(TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4_read_add),
.proj1in(TPROJ_FromPlus_F2D5_F3F4_PRD_F2D5_F3F4),
.number_in_proj2in(TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4_number),
.read_add_proj2in(TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4_read_add),
.proj2in(TPROJ_FromMinus_F2D5_F3F4_PRD_F2D5_F3F4),
.number_in_proj3in(TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4_number),
.read_add_proj3in(TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4_read_add),
.proj3in(TPROJ_F3D5F4D5_F2D5_PRD_F2D5_F3F4),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X1),
.vmprojoutPHI1X2(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X2),
.vmprojoutPHI2X1(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X1),
.vmprojoutPHI2X2(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X2),
.vmprojoutPHI3X1(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X1),
.vmprojoutPHI3X2(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X2),
.allprojout(PRD_F2D5_F3F4_AP_F3F4_F2D5),
.valid_data(PRD_F2D5_F3F4_AP_F3F4_F2D5_wr_en),
.vmprojoutPHI1X1_wr_en(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PRD_F2D5_F3F4_VMPROJ_F3F4_F2D5PHI3X2_wr_en),
.start(TPROJ_FromPlus_F2D5_F3F4_start),
.done(PRD_F2D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b0,1'b0) PRD_F5D5_F3F4(
.number_in_proj1in(TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4_number),
.read_add_proj1in(TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4_read_add),
.proj1in(TPROJ_FromPlus_F5D5_F3F4_PRD_F5D5_F3F4),
.number_in_proj2in(TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4_number),
.read_add_proj2in(TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4_read_add),
.proj2in(TPROJ_FromMinus_F5D5_F3F4_PRD_F5D5_F3F4),
.number_in_proj3in(TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4_number),
.read_add_proj3in(TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4_read_add),
.proj3in(TPROJ_F3D5F4D5_F5D5_PRD_F5D5_F3F4),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X1),
.vmprojoutPHI1X2(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X2),
.vmprojoutPHI2X1(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X1),
.vmprojoutPHI2X2(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X2),
.vmprojoutPHI3X1(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X1),
.vmprojoutPHI3X2(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X2),
.vmprojoutPHI4X1(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X1),
.vmprojoutPHI4X2(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X2),
.allprojout(PRD_F5D5_F3F4_AP_F3F4_F5D5),
.valid_data(PRD_F5D5_F3F4_AP_F3F4_F5D5_wr_en),
.vmprojoutPHI1X1_wr_en(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PRD_F5D5_F3F4_VMPROJ_F3F4_F5D5PHI4X2_wr_en),
.start(TPROJ_FromPlus_F5D5_F3F4_start),
.done(PRD_F5D5_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F3D5PHI1X1(
.number_in_vmstubin(VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1_number),
.read_add_vmstubin(VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1_read_add),
.vmstubin(VMS_F3D5PHI1X1n3_ME_F1F2_F3D5PHI1X1),
.number_in_vmprojin(VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1_read_add),
.vmprojin(VMPROJ_F1F2_F3D5PHI1X1_ME_F1F2_F3D5PHI1X1),
.matchout(ME_F1F2_F3D5PHI1X1_CM_F1F2_F3D5PHI1X1),
.valid_data(ME_F1F2_F3D5PHI1X1_CM_F1F2_F3D5PHI1X1_wr_en),
.start(VMPROJ_F1F2_F3D5PHI1X1_start),
.done(ME_F1F2_F3D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F3D5PHI1X2(
.number_in_vmstubin(VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2_number),
.read_add_vmstubin(VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2_read_add),
.vmstubin(VMS_F3D5PHI1X2n2_ME_F1F2_F3D5PHI1X2),
.number_in_vmprojin(VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2_read_add),
.vmprojin(VMPROJ_F1F2_F3D5PHI1X2_ME_F1F2_F3D5PHI1X2),
.matchout(ME_F1F2_F3D5PHI1X2_CM_F1F2_F3D5PHI1X2),
.valid_data(ME_F1F2_F3D5PHI1X2_CM_F1F2_F3D5PHI1X2_wr_en),
.start(VMPROJ_F1F2_F3D5PHI1X2_start),
.done(ME_F1F2_F3D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F3D5PHI2X1(
.number_in_vmstubin(VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1_number),
.read_add_vmstubin(VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1_read_add),
.vmstubin(VMS_F3D5PHI2X1n5_ME_F1F2_F3D5PHI2X1),
.number_in_vmprojin(VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1_read_add),
.vmprojin(VMPROJ_F1F2_F3D5PHI2X1_ME_F1F2_F3D5PHI2X1),
.matchout(ME_F1F2_F3D5PHI2X1_CM_F1F2_F3D5PHI2X1),
.valid_data(ME_F1F2_F3D5PHI2X1_CM_F1F2_F3D5PHI2X1_wr_en),
.start(VMPROJ_F1F2_F3D5PHI2X1_start),
.done(ME_F1F2_F3D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F3D5PHI2X2(
.number_in_vmstubin(VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2_number),
.read_add_vmstubin(VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2_read_add),
.vmstubin(VMS_F3D5PHI2X2n3_ME_F1F2_F3D5PHI2X2),
.number_in_vmprojin(VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2_read_add),
.vmprojin(VMPROJ_F1F2_F3D5PHI2X2_ME_F1F2_F3D5PHI2X2),
.matchout(ME_F1F2_F3D5PHI2X2_CM_F1F2_F3D5PHI2X2),
.valid_data(ME_F1F2_F3D5PHI2X2_CM_F1F2_F3D5PHI2X2_wr_en),
.start(VMPROJ_F1F2_F3D5PHI2X2_start),
.done(ME_F1F2_F3D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F3D5PHI3X1(
.number_in_vmstubin(VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1_number),
.read_add_vmstubin(VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1_read_add),
.vmstubin(VMS_F3D5PHI3X1n5_ME_F1F2_F3D5PHI3X1),
.number_in_vmprojin(VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1_read_add),
.vmprojin(VMPROJ_F1F2_F3D5PHI3X1_ME_F1F2_F3D5PHI3X1),
.matchout(ME_F1F2_F3D5PHI3X1_CM_F1F2_F3D5PHI3X1),
.valid_data(ME_F1F2_F3D5PHI3X1_CM_F1F2_F3D5PHI3X1_wr_en),
.start(VMPROJ_F1F2_F3D5PHI3X1_start),
.done(ME_F1F2_F3D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F3D5PHI3X2(
.number_in_vmstubin(VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2_number),
.read_add_vmstubin(VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2_read_add),
.vmstubin(VMS_F3D5PHI3X2n3_ME_F1F2_F3D5PHI3X2),
.number_in_vmprojin(VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2_read_add),
.vmprojin(VMPROJ_F1F2_F3D5PHI3X2_ME_F1F2_F3D5PHI3X2),
.matchout(ME_F1F2_F3D5PHI3X2_CM_F1F2_F3D5PHI3X2),
.valid_data(ME_F1F2_F3D5PHI3X2_CM_F1F2_F3D5PHI3X2_wr_en),
.start(VMPROJ_F1F2_F3D5PHI3X2_start),
.done(ME_F1F2_F3D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F3D5PHI4X1(
.number_in_vmstubin(VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1_number),
.read_add_vmstubin(VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1_read_add),
.vmstubin(VMS_F3D5PHI4X1n3_ME_F1F2_F3D5PHI4X1),
.number_in_vmprojin(VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1_read_add),
.vmprojin(VMPROJ_F1F2_F3D5PHI4X1_ME_F1F2_F3D5PHI4X1),
.matchout(ME_F1F2_F3D5PHI4X1_CM_F1F2_F3D5PHI4X1),
.valid_data(ME_F1F2_F3D5PHI4X1_CM_F1F2_F3D5PHI4X1_wr_en),
.start(VMPROJ_F1F2_F3D5PHI4X1_start),
.done(ME_F1F2_F3D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F3D5PHI4X2(
.number_in_vmstubin(VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2_number),
.read_add_vmstubin(VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2_read_add),
.vmstubin(VMS_F3D5PHI4X2n2_ME_F1F2_F3D5PHI4X2),
.number_in_vmprojin(VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2_read_add),
.vmprojin(VMPROJ_F1F2_F3D5PHI4X2_ME_F1F2_F3D5PHI4X2),
.matchout(ME_F1F2_F3D5PHI4X2_CM_F1F2_F3D5PHI4X2),
.valid_data(ME_F1F2_F3D5PHI4X2_CM_F1F2_F3D5PHI4X2_wr_en),
.start(VMPROJ_F1F2_F3D5PHI4X2_start),
.done(ME_F1F2_F3D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F4D5PHI1X1(
.number_in_vmstubin(VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1_number),
.read_add_vmstubin(VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1_read_add),
.vmstubin(VMS_F4D5PHI1X1n3_ME_F1F2_F4D5PHI1X1),
.number_in_vmprojin(VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1_read_add),
.vmprojin(VMPROJ_F1F2_F4D5PHI1X1_ME_F1F2_F4D5PHI1X1),
.matchout(ME_F1F2_F4D5PHI1X1_CM_F1F2_F4D5PHI1X1),
.valid_data(ME_F1F2_F4D5PHI1X1_CM_F1F2_F4D5PHI1X1_wr_en),
.start(VMPROJ_F1F2_F4D5PHI1X1_start),
.done(ME_F1F2_F4D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F4D5PHI1X2(
.number_in_vmstubin(VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2_number),
.read_add_vmstubin(VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2_read_add),
.vmstubin(VMS_F4D5PHI1X2n5_ME_F1F2_F4D5PHI1X2),
.number_in_vmprojin(VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2_read_add),
.vmprojin(VMPROJ_F1F2_F4D5PHI1X2_ME_F1F2_F4D5PHI1X2),
.matchout(ME_F1F2_F4D5PHI1X2_CM_F1F2_F4D5PHI1X2),
.valid_data(ME_F1F2_F4D5PHI1X2_CM_F1F2_F4D5PHI1X2_wr_en),
.start(VMPROJ_F1F2_F4D5PHI1X2_start),
.done(ME_F1F2_F4D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F4D5PHI2X1(
.number_in_vmstubin(VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1_number),
.read_add_vmstubin(VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1_read_add),
.vmstubin(VMS_F4D5PHI2X1n3_ME_F1F2_F4D5PHI2X1),
.number_in_vmprojin(VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1_read_add),
.vmprojin(VMPROJ_F1F2_F4D5PHI2X1_ME_F1F2_F4D5PHI2X1),
.matchout(ME_F1F2_F4D5PHI2X1_CM_F1F2_F4D5PHI2X1),
.valid_data(ME_F1F2_F4D5PHI2X1_CM_F1F2_F4D5PHI2X1_wr_en),
.start(VMPROJ_F1F2_F4D5PHI2X1_start),
.done(ME_F1F2_F4D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F4D5PHI2X2(
.number_in_vmstubin(VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2_number),
.read_add_vmstubin(VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2_read_add),
.vmstubin(VMS_F4D5PHI2X2n5_ME_F1F2_F4D5PHI2X2),
.number_in_vmprojin(VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2_read_add),
.vmprojin(VMPROJ_F1F2_F4D5PHI2X2_ME_F1F2_F4D5PHI2X2),
.matchout(ME_F1F2_F4D5PHI2X2_CM_F1F2_F4D5PHI2X2),
.valid_data(ME_F1F2_F4D5PHI2X2_CM_F1F2_F4D5PHI2X2_wr_en),
.start(VMPROJ_F1F2_F4D5PHI2X2_start),
.done(ME_F1F2_F4D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F4D5PHI3X1(
.number_in_vmstubin(VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1_number),
.read_add_vmstubin(VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1_read_add),
.vmstubin(VMS_F4D5PHI3X1n3_ME_F1F2_F4D5PHI3X1),
.number_in_vmprojin(VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1_read_add),
.vmprojin(VMPROJ_F1F2_F4D5PHI3X1_ME_F1F2_F4D5PHI3X1),
.matchout(ME_F1F2_F4D5PHI3X1_CM_F1F2_F4D5PHI3X1),
.valid_data(ME_F1F2_F4D5PHI3X1_CM_F1F2_F4D5PHI3X1_wr_en),
.start(VMPROJ_F1F2_F4D5PHI3X1_start),
.done(ME_F1F2_F4D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F4D5PHI3X2(
.number_in_vmstubin(VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2_number),
.read_add_vmstubin(VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2_read_add),
.vmstubin(VMS_F4D5PHI3X2n5_ME_F1F2_F4D5PHI3X2),
.number_in_vmprojin(VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2_read_add),
.vmprojin(VMPROJ_F1F2_F4D5PHI3X2_ME_F1F2_F4D5PHI3X2),
.matchout(ME_F1F2_F4D5PHI3X2_CM_F1F2_F4D5PHI3X2),
.valid_data(ME_F1F2_F4D5PHI3X2_CM_F1F2_F4D5PHI3X2_wr_en),
.start(VMPROJ_F1F2_F4D5PHI3X2_start),
.done(ME_F1F2_F4D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F5D5PHI1X1(
.number_in_vmprojin(VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1_read_add),
.vmprojin(VMPROJ_F1F2_F5D5PHI1X1_ME_F1F2_F5D5PHI1X1),
.number_in_vmstubin(VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1_number),
.read_add_vmstubin(VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1_read_add),
.vmstubin(VMS_F5D5PHI1X1n1_ME_F1F2_F5D5PHI1X1),
.matchout(ME_F1F2_F5D5PHI1X1_CM_F1F2_F5D5PHI1X1),
.valid_data(ME_F1F2_F5D5PHI1X1_CM_F1F2_F5D5PHI1X1_wr_en),
.start(VMPROJ_F1F2_F5D5PHI1X1_start),
.done(ME_F1F2_F5D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F5D5PHI1X2(
.number_in_vmprojin(VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2_read_add),
.vmprojin(VMPROJ_F1F2_F5D5PHI1X2_ME_F1F2_F5D5PHI1X2),
.number_in_vmstubin(VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2_number),
.read_add_vmstubin(VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2_read_add),
.vmstubin(VMS_F5D5PHI1X2n1_ME_F1F2_F5D5PHI1X2),
.matchout(ME_F1F2_F5D5PHI1X2_CM_F1F2_F5D5PHI1X2),
.valid_data(ME_F1F2_F5D5PHI1X2_CM_F1F2_F5D5PHI1X2_wr_en),
.start(VMPROJ_F1F2_F5D5PHI1X2_start),
.done(ME_F1F2_F5D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F5D5PHI2X1(
.number_in_vmprojin(VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1_read_add),
.vmprojin(VMPROJ_F1F2_F5D5PHI2X1_ME_F1F2_F5D5PHI2X1),
.number_in_vmstubin(VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1_number),
.read_add_vmstubin(VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1_read_add),
.vmstubin(VMS_F5D5PHI2X1n1_ME_F1F2_F5D5PHI2X1),
.matchout(ME_F1F2_F5D5PHI2X1_CM_F1F2_F5D5PHI2X1),
.valid_data(ME_F1F2_F5D5PHI2X1_CM_F1F2_F5D5PHI2X1_wr_en),
.start(VMPROJ_F1F2_F5D5PHI2X1_start),
.done(ME_F1F2_F5D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F5D5PHI2X2(
.number_in_vmprojin(VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2_read_add),
.vmprojin(VMPROJ_F1F2_F5D5PHI2X2_ME_F1F2_F5D5PHI2X2),
.number_in_vmstubin(VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2_number),
.read_add_vmstubin(VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2_read_add),
.vmstubin(VMS_F5D5PHI2X2n1_ME_F1F2_F5D5PHI2X2),
.matchout(ME_F1F2_F5D5PHI2X2_CM_F1F2_F5D5PHI2X2),
.valid_data(ME_F1F2_F5D5PHI2X2_CM_F1F2_F5D5PHI2X2_wr_en),
.start(VMPROJ_F1F2_F5D5PHI2X2_start),
.done(ME_F1F2_F5D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F5D5PHI3X1(
.number_in_vmprojin(VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1_read_add),
.vmprojin(VMPROJ_F1F2_F5D5PHI3X1_ME_F1F2_F5D5PHI3X1),
.number_in_vmstubin(VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1_number),
.read_add_vmstubin(VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1_read_add),
.vmstubin(VMS_F5D5PHI3X1n1_ME_F1F2_F5D5PHI3X1),
.matchout(ME_F1F2_F5D5PHI3X1_CM_F1F2_F5D5PHI3X1),
.valid_data(ME_F1F2_F5D5PHI3X1_CM_F1F2_F5D5PHI3X1_wr_en),
.start(VMPROJ_F1F2_F5D5PHI3X1_start),
.done(ME_F1F2_F5D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F5D5PHI3X2(
.number_in_vmprojin(VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2_read_add),
.vmprojin(VMPROJ_F1F2_F5D5PHI3X2_ME_F1F2_F5D5PHI3X2),
.number_in_vmstubin(VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2_number),
.read_add_vmstubin(VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2_read_add),
.vmstubin(VMS_F5D5PHI3X2n1_ME_F1F2_F5D5PHI3X2),
.matchout(ME_F1F2_F5D5PHI3X2_CM_F1F2_F5D5PHI3X2),
.valid_data(ME_F1F2_F5D5PHI3X2_CM_F1F2_F5D5PHI3X2_wr_en),
.start(VMPROJ_F1F2_F5D5PHI3X2_start),
.done(ME_F1F2_F5D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F5D5PHI4X1(
.number_in_vmprojin(VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1_number),
.read_add_vmprojin(VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1_read_add),
.vmprojin(VMPROJ_F1F2_F5D5PHI4X1_ME_F1F2_F5D5PHI4X1),
.number_in_vmstubin(VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1_number),
.read_add_vmstubin(VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1_read_add),
.vmstubin(VMS_F5D5PHI4X1n1_ME_F1F2_F5D5PHI4X1),
.matchout(ME_F1F2_F5D5PHI4X1_CM_F1F2_F5D5PHI4X1),
.valid_data(ME_F1F2_F5D5PHI4X1_CM_F1F2_F5D5PHI4X1_wr_en),
.start(VMPROJ_F1F2_F5D5PHI4X1_start),
.done(ME_F1F2_F5D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F1F2_F5D5PHI4X2(
.number_in_vmprojin(VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2_number),
.read_add_vmprojin(VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2_read_add),
.vmprojin(VMPROJ_F1F2_F5D5PHI4X2_ME_F1F2_F5D5PHI4X2),
.number_in_vmstubin(VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2_number),
.read_add_vmstubin(VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2_read_add),
.vmstubin(VMS_F5D5PHI4X2n1_ME_F1F2_F5D5PHI4X2),
.matchout(ME_F1F2_F5D5PHI4X2_CM_F1F2_F5D5PHI4X2),
.valid_data(ME_F1F2_F5D5PHI4X2_CM_F1F2_F5D5PHI4X2_wr_en),
.start(VMPROJ_F1F2_F5D5PHI4X2_start),
.done(ME_F1F2_F5D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F1D5PHI1X1(
.number_in_vmstubin(VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1_number),
.read_add_vmstubin(VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1_read_add),
.vmstubin(VMS_F1D5PHI1X1n3_ME_F3F4_F1D5PHI1X1),
.number_in_vmprojin(VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1_read_add),
.vmprojin(VMPROJ_F3F4_F1D5PHI1X1_ME_F3F4_F1D5PHI1X1),
.matchout(ME_F3F4_F1D5PHI1X1_CM_F3F4_F1D5PHI1X1),
.valid_data(ME_F3F4_F1D5PHI1X1_CM_F3F4_F1D5PHI1X1_wr_en),
.start(VMPROJ_F3F4_F1D5PHI1X1_start),
.done(ME_F3F4_F1D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F1D5PHI1X2(
.number_in_vmstubin(VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2_number),
.read_add_vmstubin(VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2_read_add),
.vmstubin(VMS_F1D5PHI1X2n2_ME_F3F4_F1D5PHI1X2),
.number_in_vmprojin(VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2_read_add),
.vmprojin(VMPROJ_F3F4_F1D5PHI1X2_ME_F3F4_F1D5PHI1X2),
.matchout(ME_F3F4_F1D5PHI1X2_CM_F3F4_F1D5PHI1X2),
.valid_data(ME_F3F4_F1D5PHI1X2_CM_F3F4_F1D5PHI1X2_wr_en),
.start(VMPROJ_F3F4_F1D5PHI1X2_start),
.done(ME_F3F4_F1D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F1D5PHI2X1(
.number_in_vmstubin(VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1_number),
.read_add_vmstubin(VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1_read_add),
.vmstubin(VMS_F1D5PHI2X1n5_ME_F3F4_F1D5PHI2X1),
.number_in_vmprojin(VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1_read_add),
.vmprojin(VMPROJ_F3F4_F1D5PHI2X1_ME_F3F4_F1D5PHI2X1),
.matchout(ME_F3F4_F1D5PHI2X1_CM_F3F4_F1D5PHI2X1),
.valid_data(ME_F3F4_F1D5PHI2X1_CM_F3F4_F1D5PHI2X1_wr_en),
.start(VMPROJ_F3F4_F1D5PHI2X1_start),
.done(ME_F3F4_F1D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F1D5PHI2X2(
.number_in_vmstubin(VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2_number),
.read_add_vmstubin(VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2_read_add),
.vmstubin(VMS_F1D5PHI2X2n3_ME_F3F4_F1D5PHI2X2),
.number_in_vmprojin(VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2_read_add),
.vmprojin(VMPROJ_F3F4_F1D5PHI2X2_ME_F3F4_F1D5PHI2X2),
.matchout(ME_F3F4_F1D5PHI2X2_CM_F3F4_F1D5PHI2X2),
.valid_data(ME_F3F4_F1D5PHI2X2_CM_F3F4_F1D5PHI2X2_wr_en),
.start(VMPROJ_F3F4_F1D5PHI2X2_start),
.done(ME_F3F4_F1D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F1D5PHI3X1(
.number_in_vmstubin(VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1_number),
.read_add_vmstubin(VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1_read_add),
.vmstubin(VMS_F1D5PHI3X1n5_ME_F3F4_F1D5PHI3X1),
.number_in_vmprojin(VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1_read_add),
.vmprojin(VMPROJ_F3F4_F1D5PHI3X1_ME_F3F4_F1D5PHI3X1),
.matchout(ME_F3F4_F1D5PHI3X1_CM_F3F4_F1D5PHI3X1),
.valid_data(ME_F3F4_F1D5PHI3X1_CM_F3F4_F1D5PHI3X1_wr_en),
.start(VMPROJ_F3F4_F1D5PHI3X1_start),
.done(ME_F3F4_F1D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F1D5PHI3X2(
.number_in_vmstubin(VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2_number),
.read_add_vmstubin(VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2_read_add),
.vmstubin(VMS_F1D5PHI3X2n3_ME_F3F4_F1D5PHI3X2),
.number_in_vmprojin(VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2_read_add),
.vmprojin(VMPROJ_F3F4_F1D5PHI3X2_ME_F3F4_F1D5PHI3X2),
.matchout(ME_F3F4_F1D5PHI3X2_CM_F3F4_F1D5PHI3X2),
.valid_data(ME_F3F4_F1D5PHI3X2_CM_F3F4_F1D5PHI3X2_wr_en),
.start(VMPROJ_F3F4_F1D5PHI3X2_start),
.done(ME_F3F4_F1D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F1D5PHI4X1(
.number_in_vmstubin(VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1_number),
.read_add_vmstubin(VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1_read_add),
.vmstubin(VMS_F1D5PHI4X1n3_ME_F3F4_F1D5PHI4X1),
.number_in_vmprojin(VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1_read_add),
.vmprojin(VMPROJ_F3F4_F1D5PHI4X1_ME_F3F4_F1D5PHI4X1),
.matchout(ME_F3F4_F1D5PHI4X1_CM_F3F4_F1D5PHI4X1),
.valid_data(ME_F3F4_F1D5PHI4X1_CM_F3F4_F1D5PHI4X1_wr_en),
.start(VMPROJ_F3F4_F1D5PHI4X1_start),
.done(ME_F3F4_F1D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F1D5PHI4X2(
.number_in_vmstubin(VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2_number),
.read_add_vmstubin(VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2_read_add),
.vmstubin(VMS_F1D5PHI4X2n2_ME_F3F4_F1D5PHI4X2),
.number_in_vmprojin(VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2_read_add),
.vmprojin(VMPROJ_F3F4_F1D5PHI4X2_ME_F3F4_F1D5PHI4X2),
.matchout(ME_F3F4_F1D5PHI4X2_CM_F3F4_F1D5PHI4X2),
.valid_data(ME_F3F4_F1D5PHI4X2_CM_F3F4_F1D5PHI4X2_wr_en),
.start(VMPROJ_F3F4_F1D5PHI4X2_start),
.done(ME_F3F4_F1D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F2D5PHI1X1(
.number_in_vmstubin(VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1_number),
.read_add_vmstubin(VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1_read_add),
.vmstubin(VMS_F2D5PHI1X1n3_ME_F3F4_F2D5PHI1X1),
.number_in_vmprojin(VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1_read_add),
.vmprojin(VMPROJ_F3F4_F2D5PHI1X1_ME_F3F4_F2D5PHI1X1),
.matchout(ME_F3F4_F2D5PHI1X1_CM_F3F4_F2D5PHI1X1),
.valid_data(ME_F3F4_F2D5PHI1X1_CM_F3F4_F2D5PHI1X1_wr_en),
.start(VMPROJ_F3F4_F2D5PHI1X1_start),
.done(ME_F3F4_F2D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F2D5PHI1X2(
.number_in_vmstubin(VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2_number),
.read_add_vmstubin(VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2_read_add),
.vmstubin(VMS_F2D5PHI1X2n5_ME_F3F4_F2D5PHI1X2),
.number_in_vmprojin(VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2_read_add),
.vmprojin(VMPROJ_F3F4_F2D5PHI1X2_ME_F3F4_F2D5PHI1X2),
.matchout(ME_F3F4_F2D5PHI1X2_CM_F3F4_F2D5PHI1X2),
.valid_data(ME_F3F4_F2D5PHI1X2_CM_F3F4_F2D5PHI1X2_wr_en),
.start(VMPROJ_F3F4_F2D5PHI1X2_start),
.done(ME_F3F4_F2D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F2D5PHI2X1(
.number_in_vmstubin(VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1_number),
.read_add_vmstubin(VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1_read_add),
.vmstubin(VMS_F2D5PHI2X1n3_ME_F3F4_F2D5PHI2X1),
.number_in_vmprojin(VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1_read_add),
.vmprojin(VMPROJ_F3F4_F2D5PHI2X1_ME_F3F4_F2D5PHI2X1),
.matchout(ME_F3F4_F2D5PHI2X1_CM_F3F4_F2D5PHI2X1),
.valid_data(ME_F3F4_F2D5PHI2X1_CM_F3F4_F2D5PHI2X1_wr_en),
.start(VMPROJ_F3F4_F2D5PHI2X1_start),
.done(ME_F3F4_F2D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F2D5PHI2X2(
.number_in_vmstubin(VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2_number),
.read_add_vmstubin(VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2_read_add),
.vmstubin(VMS_F2D5PHI2X2n5_ME_F3F4_F2D5PHI2X2),
.number_in_vmprojin(VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2_read_add),
.vmprojin(VMPROJ_F3F4_F2D5PHI2X2_ME_F3F4_F2D5PHI2X2),
.matchout(ME_F3F4_F2D5PHI2X2_CM_F3F4_F2D5PHI2X2),
.valid_data(ME_F3F4_F2D5PHI2X2_CM_F3F4_F2D5PHI2X2_wr_en),
.start(VMPROJ_F3F4_F2D5PHI2X2_start),
.done(ME_F3F4_F2D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F2D5PHI3X1(
.number_in_vmstubin(VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1_number),
.read_add_vmstubin(VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1_read_add),
.vmstubin(VMS_F2D5PHI3X1n3_ME_F3F4_F2D5PHI3X1),
.number_in_vmprojin(VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1_read_add),
.vmprojin(VMPROJ_F3F4_F2D5PHI3X1_ME_F3F4_F2D5PHI3X1),
.matchout(ME_F3F4_F2D5PHI3X1_CM_F3F4_F2D5PHI3X1),
.valid_data(ME_F3F4_F2D5PHI3X1_CM_F3F4_F2D5PHI3X1_wr_en),
.start(VMPROJ_F3F4_F2D5PHI3X1_start),
.done(ME_F3F4_F2D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F2D5PHI3X2(
.number_in_vmstubin(VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2_number),
.read_add_vmstubin(VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2_read_add),
.vmstubin(VMS_F2D5PHI3X2n5_ME_F3F4_F2D5PHI3X2),
.number_in_vmprojin(VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2_read_add),
.vmprojin(VMPROJ_F3F4_F2D5PHI3X2_ME_F3F4_F2D5PHI3X2),
.matchout(ME_F3F4_F2D5PHI3X2_CM_F3F4_F2D5PHI3X2),
.valid_data(ME_F3F4_F2D5PHI3X2_CM_F3F4_F2D5PHI3X2_wr_en),
.start(VMPROJ_F3F4_F2D5PHI3X2_start),
.done(ME_F3F4_F2D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F5D5PHI1X1(
.number_in_vmstubin(VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1_number),
.read_add_vmstubin(VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1_read_add),
.vmstubin(VMS_F5D5PHI1X1n2_ME_F3F4_F5D5PHI1X1),
.number_in_vmprojin(VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1_read_add),
.vmprojin(VMPROJ_F3F4_F5D5PHI1X1_ME_F3F4_F5D5PHI1X1),
.matchout(ME_F3F4_F5D5PHI1X1_CM_F3F4_F5D5PHI1X1),
.valid_data(ME_F3F4_F5D5PHI1X1_CM_F3F4_F5D5PHI1X1_wr_en),
.start(VMPROJ_F3F4_F5D5PHI1X1_start),
.done(ME_F3F4_F5D5PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F5D5PHI1X2(
.number_in_vmstubin(VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2_number),
.read_add_vmstubin(VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2_read_add),
.vmstubin(VMS_F5D5PHI1X2n2_ME_F3F4_F5D5PHI1X2),
.number_in_vmprojin(VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2_read_add),
.vmprojin(VMPROJ_F3F4_F5D5PHI1X2_ME_F3F4_F5D5PHI1X2),
.matchout(ME_F3F4_F5D5PHI1X2_CM_F3F4_F5D5PHI1X2),
.valid_data(ME_F3F4_F5D5PHI1X2_CM_F3F4_F5D5PHI1X2_wr_en),
.start(VMPROJ_F3F4_F5D5PHI1X2_start),
.done(ME_F3F4_F5D5PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F5D5PHI2X1(
.number_in_vmstubin(VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1_number),
.read_add_vmstubin(VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1_read_add),
.vmstubin(VMS_F5D5PHI2X1n2_ME_F3F4_F5D5PHI2X1),
.number_in_vmprojin(VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1_read_add),
.vmprojin(VMPROJ_F3F4_F5D5PHI2X1_ME_F3F4_F5D5PHI2X1),
.matchout(ME_F3F4_F5D5PHI2X1_CM_F3F4_F5D5PHI2X1),
.valid_data(ME_F3F4_F5D5PHI2X1_CM_F3F4_F5D5PHI2X1_wr_en),
.start(VMPROJ_F3F4_F5D5PHI2X1_start),
.done(ME_F3F4_F5D5PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F5D5PHI2X2(
.number_in_vmstubin(VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2_number),
.read_add_vmstubin(VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2_read_add),
.vmstubin(VMS_F5D5PHI2X2n2_ME_F3F4_F5D5PHI2X2),
.number_in_vmprojin(VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2_read_add),
.vmprojin(VMPROJ_F3F4_F5D5PHI2X2_ME_F3F4_F5D5PHI2X2),
.matchout(ME_F3F4_F5D5PHI2X2_CM_F3F4_F5D5PHI2X2),
.valid_data(ME_F3F4_F5D5PHI2X2_CM_F3F4_F5D5PHI2X2_wr_en),
.start(VMPROJ_F3F4_F5D5PHI2X2_start),
.done(ME_F3F4_F5D5PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F5D5PHI3X1(
.number_in_vmstubin(VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1_number),
.read_add_vmstubin(VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1_read_add),
.vmstubin(VMS_F5D5PHI3X1n2_ME_F3F4_F5D5PHI3X1),
.number_in_vmprojin(VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1_read_add),
.vmprojin(VMPROJ_F3F4_F5D5PHI3X1_ME_F3F4_F5D5PHI3X1),
.matchout(ME_F3F4_F5D5PHI3X1_CM_F3F4_F5D5PHI3X1),
.valid_data(ME_F3F4_F5D5PHI3X1_CM_F3F4_F5D5PHI3X1_wr_en),
.start(VMPROJ_F3F4_F5D5PHI3X1_start),
.done(ME_F3F4_F5D5PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F5D5PHI3X2(
.number_in_vmstubin(VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2_number),
.read_add_vmstubin(VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2_read_add),
.vmstubin(VMS_F5D5PHI3X2n2_ME_F3F4_F5D5PHI3X2),
.number_in_vmprojin(VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2_read_add),
.vmprojin(VMPROJ_F3F4_F5D5PHI3X2_ME_F3F4_F5D5PHI3X2),
.matchout(ME_F3F4_F5D5PHI3X2_CM_F3F4_F5D5PHI3X2),
.valid_data(ME_F3F4_F5D5PHI3X2_CM_F3F4_F5D5PHI3X2_wr_en),
.start(VMPROJ_F3F4_F5D5PHI3X2_start),
.done(ME_F3F4_F5D5PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F5D5PHI4X1(
.number_in_vmstubin(VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1_number),
.read_add_vmstubin(VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1_read_add),
.vmstubin(VMS_F5D5PHI4X1n2_ME_F3F4_F5D5PHI4X1),
.number_in_vmprojin(VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1_number),
.read_add_vmprojin(VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1_read_add),
.vmprojin(VMPROJ_F3F4_F5D5PHI4X1_ME_F3F4_F5D5PHI4X1),
.matchout(ME_F3F4_F5D5PHI4X1_CM_F3F4_F5D5PHI4X1),
.valid_data(ME_F3F4_F5D5PHI4X1_CM_F3F4_F5D5PHI4X1_wr_en),
.start(VMPROJ_F3F4_F5D5PHI4X1_start),
.done(ME_F3F4_F5D5PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_F3F4_F5D5PHI4X2(
.number_in_vmstubin(VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2_number),
.read_add_vmstubin(VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2_read_add),
.vmstubin(VMS_F5D5PHI4X2n2_ME_F3F4_F5D5PHI4X2),
.number_in_vmprojin(VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2_number),
.read_add_vmprojin(VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2_read_add),
.vmprojin(VMPROJ_F3F4_F5D5PHI4X2_ME_F3F4_F5D5PHI4X2),
.matchout(ME_F3F4_F5D5PHI4X2_CM_F3F4_F5D5PHI4X2),
.valid_data(ME_F3F4_F5D5PHI4X2_CM_F3F4_F5D5PHI4X2_wr_en),
.start(VMPROJ_F3F4_F5D5PHI4X2_start),
.done(ME_F3F4_F5D5PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

DiskMatchCalculator #(3'b100,1'b1) MC_F1F2_F3D5(
.number_in_match1in(CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5_number),
.read_add_match1in(CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5_read_add),
.match1in(CM_F1F2_F3D5PHI1X1_MC_F1F2_F3D5),
.number_in_match2in(CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5_number),
.read_add_match2in(CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5_read_add),
.match2in(CM_F1F2_F3D5PHI1X2_MC_F1F2_F3D5),
.number_in_match3in(CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5_number),
.read_add_match3in(CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5_read_add),
.match3in(CM_F1F2_F3D5PHI2X1_MC_F1F2_F3D5),
.number_in_match4in(CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5_number),
.read_add_match4in(CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5_read_add),
.match4in(CM_F1F2_F3D5PHI2X2_MC_F1F2_F3D5),
.number_in_match5in(CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5_number),
.read_add_match5in(CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5_read_add),
.match5in(CM_F1F2_F3D5PHI3X1_MC_F1F2_F3D5),
.number_in_match6in(CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5_number),
.read_add_match6in(CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5_read_add),
.match6in(CM_F1F2_F3D5PHI3X2_MC_F1F2_F3D5),
.number_in_match7in(CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5_number),
.read_add_match7in(CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5_read_add),
.match7in(CM_F1F2_F3D5PHI4X1_MC_F1F2_F3D5),
.number_in_match8in(CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5_number),
.read_add_match8in(CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5_read_add),
.match8in(CM_F1F2_F3D5PHI4X2_MC_F1F2_F3D5),
.read_add_allprojin(AP_F1F2_F3D5_MC_F1F2_F3D5_read_add),
.allprojin(AP_F1F2_F3D5_MC_F1F2_F3D5),
.read_add_allstubin(AS_F3D5n2_MC_F1F2_F3D5_read_add),
.allstubin(AS_F3D5n2_MC_F1F2_F3D5),
.matchoutminus(MC_F1F2_F3D5_FM_F1F2_F3D5_ToMinus),
.matchoutplus(MC_F1F2_F3D5_FM_F1F2_F3D5_ToPlus),
.matchout1(MC_F1F2_F3D5_FM_F1F2_F3D5),
.valid_matchminus(MC_F1F2_F3D5_FM_F1F2_F3D5_ToMinus_wr_en),
.valid_matchplus(MC_F1F2_F3D5_FM_F1F2_F3D5_ToPlus_wr_en),
.valid_match(MC_F1F2_F3D5_FM_F1F2_F3D5_wr_en),
.start(CM_F1F2_F3D5PHI1X1_start),
.done(MC_F1F2_F3D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

DiskMatchCalculator #(3'b100,1'b1) MC_F1F2_F4D5(
.number_in_match1in(CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5_number),
.read_add_match1in(CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5_read_add),
.match1in(CM_F1F2_F4D5PHI1X1_MC_F1F2_F4D5),
.number_in_match2in(CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5_number),
.read_add_match2in(CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5_read_add),
.match2in(CM_F1F2_F4D5PHI1X2_MC_F1F2_F4D5),
.number_in_match3in(CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5_number),
.read_add_match3in(CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5_read_add),
.match3in(CM_F1F2_F4D5PHI2X1_MC_F1F2_F4D5),
.number_in_match4in(CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5_number),
.read_add_match4in(CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5_read_add),
.match4in(CM_F1F2_F4D5PHI2X2_MC_F1F2_F4D5),
.number_in_match5in(CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5_number),
.read_add_match5in(CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5_read_add),
.match5in(CM_F1F2_F4D5PHI3X1_MC_F1F2_F4D5),
.number_in_match6in(CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5_number),
.read_add_match6in(CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5_read_add),
.match6in(CM_F1F2_F4D5PHI3X2_MC_F1F2_F4D5),
.read_add_allprojin(AP_F1F2_F4D5_MC_F1F2_F4D5_read_add),
.allprojin(AP_F1F2_F4D5_MC_F1F2_F4D5),
.read_add_allstubin(AS_F4D5n2_MC_F1F2_F4D5_read_add),
.allstubin(AS_F4D5n2_MC_F1F2_F4D5),
.matchoutminus(MC_F1F2_F4D5_FM_F1F2_F4D5_ToMinus),
.matchoutplus(MC_F1F2_F4D5_FM_F1F2_F4D5_ToPlus),
.matchout1(MC_F1F2_F4D5_FM_F1F2_F4D5),
.valid_matchminus(MC_F1F2_F4D5_FM_F1F2_F4D5_ToMinus_wr_en),
.valid_matchplus(MC_F1F2_F4D5_FM_F1F2_F4D5_ToPlus_wr_en),
.valid_match(MC_F1F2_F4D5_FM_F1F2_F4D5_wr_en),
.start(CM_F1F2_F4D5PHI1X1_start),
.done(MC_F1F2_F4D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

DiskMatchCalculator #(3'b100,1'b1) MC_F1F2_F5D5(
.number_in_match1in(CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5_number),
.read_add_match1in(CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5_read_add),
.match1in(CM_F1F2_F5D5PHI1X1_MC_F1F2_F5D5),
.number_in_match2in(CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5_number),
.read_add_match2in(CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5_read_add),
.match2in(CM_F1F2_F5D5PHI1X2_MC_F1F2_F5D5),
.number_in_match3in(CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5_number),
.read_add_match3in(CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5_read_add),
.match3in(CM_F1F2_F5D5PHI2X1_MC_F1F2_F5D5),
.number_in_match4in(CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5_number),
.read_add_match4in(CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5_read_add),
.match4in(CM_F1F2_F5D5PHI2X2_MC_F1F2_F5D5),
.number_in_match5in(CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5_number),
.read_add_match5in(CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5_read_add),
.match5in(CM_F1F2_F5D5PHI3X1_MC_F1F2_F5D5),
.number_in_match6in(CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5_number),
.read_add_match6in(CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5_read_add),
.match6in(CM_F1F2_F5D5PHI3X2_MC_F1F2_F5D5),
.number_in_match7in(CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5_number),
.read_add_match7in(CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5_read_add),
.match7in(CM_F1F2_F5D5PHI4X1_MC_F1F2_F5D5),
.number_in_match8in(CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5_number),
.read_add_match8in(CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5_read_add),
.match8in(CM_F1F2_F5D5PHI4X2_MC_F1F2_F5D5),
.read_add_allprojin(AP_F1F2_F5D5_MC_F1F2_F5D5_read_add),
.allprojin(AP_F1F2_F5D5_MC_F1F2_F5D5),
.read_add_allstubin(AS_F5D5n1_MC_F1F2_F5D5_read_add),
.allstubin(AS_F5D5n1_MC_F1F2_F5D5),
.matchoutminus(MC_F1F2_F5D5_FM_F1F2_F5D5_ToMinus),
.matchoutplus(MC_F1F2_F5D5_FM_F1F2_F5D5_ToPlus),
.matchout1(MC_F1F2_F5D5_FM_F1F2_F5D5),
.valid_matchminus(MC_F1F2_F5D5_FM_F1F2_F5D5_ToMinus_wr_en),
.valid_matchplus(MC_F1F2_F5D5_FM_F1F2_F5D5_ToPlus_wr_en),
.valid_match(MC_F1F2_F5D5_FM_F1F2_F5D5_wr_en),
.start(CM_F1F2_F5D5PHI1X1_start),
.done(MC_F1F2_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

DiskMatchCalculator #(3'b100,1'b1) MC_F3F4_F1D5(
.number_in_match1in(CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5_number),
.read_add_match1in(CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5_read_add),
.match1in(CM_F3F4_F1D5PHI1X1_MC_F3F4_F1D5),
.number_in_match2in(CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5_number),
.read_add_match2in(CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5_read_add),
.match2in(CM_F3F4_F1D5PHI1X2_MC_F3F4_F1D5),
.number_in_match3in(CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5_number),
.read_add_match3in(CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5_read_add),
.match3in(CM_F3F4_F1D5PHI2X1_MC_F3F4_F1D5),
.number_in_match4in(CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5_number),
.read_add_match4in(CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5_read_add),
.match4in(CM_F3F4_F1D5PHI2X2_MC_F3F4_F1D5),
.number_in_match5in(CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5_number),
.read_add_match5in(CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5_read_add),
.match5in(CM_F3F4_F1D5PHI3X1_MC_F3F4_F1D5),
.number_in_match6in(CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5_number),
.read_add_match6in(CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5_read_add),
.match6in(CM_F3F4_F1D5PHI3X2_MC_F3F4_F1D5),
.number_in_match7in(CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5_number),
.read_add_match7in(CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5_read_add),
.match7in(CM_F3F4_F1D5PHI4X1_MC_F3F4_F1D5),
.number_in_match8in(CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5_number),
.read_add_match8in(CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5_read_add),
.match8in(CM_F3F4_F1D5PHI4X2_MC_F3F4_F1D5),
.read_add_allprojin(AP_F3F4_F1D5_MC_F3F4_F1D5_read_add),
.allprojin(AP_F3F4_F1D5_MC_F3F4_F1D5),
.read_add_allstubin(AS_F1D5n2_MC_F3F4_F1D5_read_add),
.allstubin(AS_F1D5n2_MC_F3F4_F1D5),
.matchoutminus(MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToMinus),
.matchoutplus(MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToPlus),
.matchout1(MC_F3F4_F1D5_FM_F3F4_F1D5),
.valid_matchminus(MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToMinus_wr_en),
.valid_matchplus(MC_F3F4_F1D5_FM_FL3FL4_F1D5_ToPlus_wr_en),
.valid_match(MC_F3F4_F1D5_FM_F3F4_F1D5_wr_en),
.start(CM_F3F4_F1D5PHI1X1_start),
.done(MC_F3F4_F1D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

DiskMatchCalculator #(3'b100,1'b1) MC_F3F4_F2D5(
.number_in_match1in(CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5_number),
.read_add_match1in(CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5_read_add),
.match1in(CM_F3F4_F2D5PHI1X1_MC_F3F4_F2D5),
.number_in_match2in(CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5_number),
.read_add_match2in(CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5_read_add),
.match2in(CM_F3F4_F2D5PHI1X2_MC_F3F4_F2D5),
.number_in_match3in(CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5_number),
.read_add_match3in(CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5_read_add),
.match3in(CM_F3F4_F2D5PHI2X1_MC_F3F4_F2D5),
.number_in_match4in(CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5_number),
.read_add_match4in(CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5_read_add),
.match4in(CM_F3F4_F2D5PHI2X2_MC_F3F4_F2D5),
.number_in_match5in(CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5_number),
.read_add_match5in(CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5_read_add),
.match5in(CM_F3F4_F2D5PHI3X1_MC_F3F4_F2D5),
.number_in_match6in(CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5_number),
.read_add_match6in(CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5_read_add),
.match6in(CM_F3F4_F2D5PHI3X2_MC_F3F4_F2D5),
.read_add_allprojin(AP_F3F4_F2D5_MC_F3F4_F2D5_read_add),
.allprojin(AP_F3F4_F2D5_MC_F3F4_F2D5),
.read_add_allstubin(AS_F2D5n2_MC_F3F4_F2D5_read_add),
.allstubin(AS_F2D5n2_MC_F3F4_F2D5),
.matchoutminus(MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToMinus),
.matchoutplus(MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToPlus),
.matchout1(MC_F3F4_F2D5_FM_F3F4_F2D5),
.valid_matchminus(MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToMinus_wr_en),
.valid_matchplus(MC_F3F4_F2D5_FM_FL3FL4_F2D5_ToPlus_wr_en),
.valid_match(MC_F3F4_F2D5_FM_F3F4_F2D5_wr_en),
.start(CM_F3F4_F2D5PHI1X1_start),
.done(MC_F3F4_F2D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

DiskMatchCalculator #(3'b100,1'b1) MC_F3F4_F5D5(
.number_in_match1in(CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5_number),
.read_add_match1in(CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5_read_add),
.match1in(CM_F3F4_F5D5PHI1X1_MC_F3F4_F5D5),
.number_in_match2in(CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5_number),
.read_add_match2in(CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5_read_add),
.match2in(CM_F3F4_F5D5PHI1X2_MC_F3F4_F5D5),
.number_in_match3in(CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5_number),
.read_add_match3in(CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5_read_add),
.match3in(CM_F3F4_F5D5PHI2X1_MC_F3F4_F5D5),
.number_in_match4in(CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5_number),
.read_add_match4in(CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5_read_add),
.match4in(CM_F3F4_F5D5PHI2X2_MC_F3F4_F5D5),
.number_in_match5in(CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5_number),
.read_add_match5in(CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5_read_add),
.match5in(CM_F3F4_F5D5PHI3X1_MC_F3F4_F5D5),
.number_in_match6in(CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5_number),
.read_add_match6in(CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5_read_add),
.match6in(CM_F3F4_F5D5PHI3X2_MC_F3F4_F5D5),
.number_in_match7in(CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5_number),
.read_add_match7in(CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5_read_add),
.match7in(CM_F3F4_F5D5PHI4X1_MC_F3F4_F5D5),
.number_in_match8in(CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5_number),
.read_add_match8in(CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5_read_add),
.match8in(CM_F3F4_F5D5PHI4X2_MC_F3F4_F5D5),
.read_add_allprojin(AP_F3F4_F5D5_MC_F3F4_F5D5_read_add),
.allprojin(AP_F3F4_F5D5_MC_F3F4_F5D5),
.read_add_allstubin(AS_F5D5n2_MC_F3F4_F5D5_read_add),
.allstubin(AS_F5D5n2_MC_F3F4_F5D5),
.matchoutminus(MC_F3F4_F5D5_FM_F3F4_F5D5_ToMinus),
.matchoutplus(MC_F3F4_F5D5_FM_F3F4_F5D5_ToPlus),
.matchout1(MC_F3F4_F5D5_FM_F3F4_F5D5),
.valid_matchminus(MC_F3F4_F5D5_FM_F3F4_F5D5_ToMinus_wr_en),
.valid_matchplus(MC_F3F4_F5D5_FM_F3F4_F5D5_ToPlus_wr_en),
.valid_match(MC_F3F4_F5D5_FM_F3F4_F5D5_wr_en),
.start(CM_F3F4_F5D5PHI1X1_start),
.done(MC_F3F4_F5D5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchTransceiver #("Disk") MT_FDSK_Minus(
.number_in_proj1in(FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus_number),
.read_add_proj1in(FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus_read_add),
.proj1in(FM_F1F2_F3D5_ToMinus_MT_FDSK_Minus),
.number_in_proj2in(FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus_number),
.read_add_proj2in(FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus_read_add),
.proj2in(FM_F1F2_F4D5_ToMinus_MT_FDSK_Minus),
.number_in_proj3in(FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus_number),
.read_add_proj3in(FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus_read_add),
.proj3in(FM_F1F2_F5D5_ToMinus_MT_FDSK_Minus),
.number_in_proj4in(FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus_number),
.read_add_proj4in(FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus_read_add),
.proj4in(FM_FL3FL4_F1D5_ToMinus_MT_FDSK_Minus),
.number_in_proj5in(FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus_number),
.read_add_proj5in(FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus_read_add),
.proj5in(FM_FL3FL4_F2D5_ToMinus_MT_FDSK_Minus),
.number_in_proj6in(FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus_number),
.read_add_proj6in(FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus_read_add),
.proj6in(FM_F3F4_F5D5_ToMinus_MT_FDSK_Minus),
.valid_incomming_match_data_stream(MT_FDSK_Minus_From_DataStream_en),
.incomming_match_data_stream(MT_FDSK_Minus_From_DataStream),
.number_in_proj7in(6'b0),
.number_in_proj8in(6'b0),
.number_in_proj9in(6'b0),
.number_in_proj10in(6'b0),
.number_in_proj11in(6'b0),
.number_in_proj12in(6'b0),
.number_in_proj13in(6'b0),
.number_in_proj14in(6'b0),
.number_in_proj15in(6'b0),
.number_in_proj16in(6'b0),
.number_in_proj17in(6'b0),
.number_in_proj18in(6'b0),
.number_in_proj19in(6'b0),
.number_in_proj20in(6'b0),
.number_in_proj21in(6'b0),
.number_in_proj22in(6'b0),
.number_in_proj23in(6'b0),
.number_in_proj24in(6'b0),
.matchout1(MT_FDSK_Minus_FM_F1F2_F3_FromMinus),
.matchout2(MT_FDSK_Minus_FM_F1F2_F4_FromMinus),
.matchout3(MT_FDSK_Minus_FM_F1F2_F5_FromMinus),
.matchout4(MT_FDSK_Minus_FM_F3F4_F1_FromMinus),
.matchout5(MT_FDSK_Minus_FM_F3F4_F2_FromMinus),
.matchout6(MT_FDSK_Minus_FM_F3F4_F5_FromMinus),
.valid_matchout1(MT_FDSK_Minus_FM_F1F2_F3_FromMinus_wr_en),
.valid_matchout2(MT_FDSK_Minus_FM_F1F2_F4_FromMinus_wr_en),
.valid_matchout3(MT_FDSK_Minus_FM_F1F2_F5_FromMinus_wr_en),
.valid_matchout4(MT_FDSK_Minus_FM_F3F4_F1_FromMinus_wr_en),
.valid_matchout5(MT_FDSK_Minus_FM_F3F4_F2_FromMinus_wr_en),
.valid_matchout6(MT_FDSK_Minus_FM_F3F4_F5_FromMinus_wr_en),
.valid_match_data_stream(MT_FDSK_Minus_To_DataStream_en),
.match_data_stream(MT_FDSK_Minus_To_DataStream),
.start(FM_F1F2_F3D5_ToMinus_start),
.done(MT_FDSK_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchTransceiver #("Disk") MT_FDSK_Plus(
.number_in_proj1in(FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus_number),
.read_add_proj1in(FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus_read_add),
.proj1in(FM_F1F2_F3D5_ToPlus_MT_FDSK_Plus),
.number_in_proj2in(FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus_number),
.read_add_proj2in(FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus_read_add),
.proj2in(FM_F1F2_F4D5_ToPlus_MT_FDSK_Plus),
.number_in_proj3in(FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus_number),
.read_add_proj3in(FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus_read_add),
.proj3in(FM_F1F2_F5D5_ToPlus_MT_FDSK_Plus),
.number_in_proj4in(FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus_number),
.read_add_proj4in(FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus_read_add),
.proj4in(FM_FL3FL4_F1D5_ToPlus_MT_FDSK_Plus),
.number_in_proj5in(FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus_number),
.read_add_proj5in(FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus_read_add),
.proj5in(FM_FL3FL4_F2D5_ToPlus_MT_FDSK_Plus),
.number_in_proj6in(FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus_number),
.read_add_proj6in(FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus_read_add),
.proj6in(FM_F3F4_F5D5_ToPlus_MT_FDSK_Plus),
.valid_incomming_match_data_stream(MT_FDSK_Plus_From_DataStream_en),
.incomming_match_data_stream(MT_FDSK_Plus_From_DataStream),
.number_in_proj7in(6'b0),
.number_in_proj8in(6'b0),
.number_in_proj9in(6'b0),
.number_in_proj10in(6'b0),
.number_in_proj11in(6'b0),
.number_in_proj12in(6'b0),
.number_in_proj13in(6'b0),
.number_in_proj14in(6'b0),
.number_in_proj15in(6'b0),
.number_in_proj16in(6'b0),
.number_in_proj17in(6'b0),
.number_in_proj18in(6'b0),
.number_in_proj19in(6'b0),
.number_in_proj20in(6'b0),
.number_in_proj21in(6'b0),
.number_in_proj22in(6'b0),
.number_in_proj23in(6'b0),
.number_in_proj24in(6'b0),
.matchout1(MT_FDSK_Plus_FM_F1F2_F3_FromPlus),
.matchout2(MT_FDSK_Plus_FM_F1F2_F4_FromPlus),
.matchout3(MT_FDSK_Plus_FM_F1F2_F5_FromPlus),
.matchout4(MT_FDSK_Plus_FM_F3F4_F1_FromPlus),
.matchout5(MT_FDSK_Plus_FM_F3F4_F2_FromPlus),
.matchout6(MT_FDSK_Plus_FM_F3F4_F5_FromPlus),
.valid_matchout1(MT_FDSK_Plus_FM_F1F2_F3_FromPlus_wr_en),
.valid_matchout2(MT_FDSK_Plus_FM_F1F2_F4_FromPlus_wr_en),
.valid_matchout3(MT_FDSK_Plus_FM_F1F2_F5_FromPlus_wr_en),
.valid_matchout4(MT_FDSK_Plus_FM_F3F4_F1_FromPlus_wr_en),
.valid_matchout5(MT_FDSK_Plus_FM_F3F4_F2_FromPlus_wr_en),
.valid_matchout6(MT_FDSK_Plus_FM_F3F4_F5_FromPlus_wr_en),
.valid_match_data_stream(MT_FDSK_Plus_To_DataStream_en),
.match_data_stream(MT_FDSK_Plus_To_DataStream),
.start(FM_F1F2_F3D5_ToPlus_start),
.done(MT_FDSK_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

FitTrack #("F1F2") FT_F1F2(
.number3in1(FM_F1F2_F3D5_FT_F1F2_number),
.read_add3in1(FM_F1F2_F3D5_FT_F1F2_read_add),
.read_en3in1(FM_F1F2_F3D5_FT_F1F2_read_en),
.fullmatch3in1(FM_F1F2_F3D5_FT_F1F2),
.number4in1(FM_F1F2_F4D5_FT_F1F2_number),
.read_add4in1(FM_F1F2_F4D5_FT_F1F2_read_add),
.read_en4in1(FM_F1F2_F4D5_FT_F1F2_read_en),
.fullmatch4in1(FM_F1F2_F4D5_FT_F1F2),
.number5in1(FM_F1F2_F5D5_FT_F1F2_number),
.read_add5in1(FM_F1F2_F5D5_FT_F1F2_read_add),
.read_en5in1(FM_F1F2_F5D5_FT_F1F2_read_en),
.fullmatch5in1(FM_F1F2_F5D5_FT_F1F2),
.read_add_pars1(TPAR_F1D5F2D5_FT_F1F2_read_add),
.tpar1in(TPAR_F1D5F2D5_FT_F1F2),
.number3in2(FM_F1F2_F3_FromMinus_FT_F1F2_number),
.read_add3in2(FM_F1F2_F3_FromMinus_FT_F1F2_read_add),
.read_en3in2(FM_F1F2_F3_FromMinus_FT_F1F2_read_en),
.fullmatch3in2(FM_F1F2_F3_FromMinus_FT_F1F2),
.number4in2(FM_F1F2_F4_FromMinus_FT_F1F2_number),
.read_add4in2(FM_F1F2_F4_FromMinus_FT_F1F2_read_add),
.read_en4in2(FM_F1F2_F4_FromMinus_FT_F1F2_read_en),
.fullmatch4in2(FM_F1F2_F4_FromMinus_FT_F1F2),
.number5in2(FM_F1F2_F5_FromMinus_FT_F1F2_number),
.read_add5in2(FM_F1F2_F5_FromMinus_FT_F1F2_read_add),
.read_en5in2(FM_F1F2_F5_FromMinus_FT_F1F2_read_en),
.fullmatch5in2(FM_F1F2_F5_FromMinus_FT_F1F2),
.number3in3(FM_F1F2_F3_FromPlus_FT_F1F2_number),
.read_add3in3(FM_F1F2_F3_FromPlus_FT_F1F2_read_add),
.read_en3in3(FM_F1F2_F3_FromPlus_FT_F1F2_read_en),
.fullmatch3in3(FM_F1F2_F3_FromPlus_FT_F1F2),
.number4in3(FM_F1F2_F4_FromPlus_FT_F1F2_number),
.read_add4in3(FM_F1F2_F4_FromPlus_FT_F1F2_read_add),
.read_en4in3(FM_F1F2_F4_FromPlus_FT_F1F2_read_en),
.fullmatch4in3(FM_F1F2_F4_FromPlus_FT_F1F2),
.number5in3(FM_F1F2_F5_FromPlus_FT_F1F2_number),
.read_add5in3(FM_F1F2_F5_FromPlus_FT_F1F2_read_add),
.read_en5in3(FM_F1F2_F5_FromPlus_FT_F1F2_read_en),
.fullmatch5in3(FM_F1F2_F5_FromPlus_FT_F1F2),
.trackout(FT_F1F2_TF_F1F2),
.valid_fit(FT_F1F2_TF_F1F2_wr_en),
.start(FM_F1F2_F5_FromPlus_start),
.done(FT_F1F2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

FitTrack #("F3F4") FT_F3F4(
.number3in1(FM_F3F4_F1D5_FT_F3F4_number),
.read_add3in1(FM_F3F4_F1D5_FT_F3F4_read_add),
.read_en3in1(FM_F3F4_F1D5_FT_F3F4_read_en),
.fullmatch3in1(FM_F3F4_F1D5_FT_F3F4),
.number4in1(FM_F3F4_F2D5_FT_F3F4_number),
.read_add4in1(FM_F3F4_F2D5_FT_F3F4_read_add),
.read_en4in1(FM_F3F4_F2D5_FT_F3F4_read_en),
.fullmatch4in1(FM_F3F4_F2D5_FT_F3F4),
.number5in1(FM_F3F4_F5D5_FT_F3F4_number),
.read_add5in1(FM_F3F4_F5D5_FT_F3F4_read_add),
.read_en5in1(FM_F3F4_F5D5_FT_F3F4_read_en),
.fullmatch5in1(FM_F3F4_F5D5_FT_F3F4),
.read_add_pars1(TPAR_F3D5F4D5_FT_F3F4_read_add),
.tpar1in(TPAR_F3D5F4D5_FT_F3F4),
.number3in2(FM_F3F4_F1_FromMinus_FT_F3F4_number),
.read_add3in2(FM_F3F4_F1_FromMinus_FT_F3F4_read_add),
.read_en3in2(FM_F3F4_F1_FromMinus_FT_F3F4_read_en),
.fullmatch3in2(FM_F3F4_F1_FromMinus_FT_F3F4),
.number4in2(FM_F3F4_F2_FromMinus_FT_F3F4_number),
.read_add4in2(FM_F3F4_F2_FromMinus_FT_F3F4_read_add),
.read_en4in2(FM_F3F4_F2_FromMinus_FT_F3F4_read_en),
.fullmatch4in2(FM_F3F4_F2_FromMinus_FT_F3F4),
.number5in2(FM_F3F4_F5_FromMinus_FT_F3F4_number),
.read_add5in2(FM_F3F4_F5_FromMinus_FT_F3F4_read_add),
.read_en5in2(FM_F3F4_F5_FromMinus_FT_F3F4_read_en),
.fullmatch5in2(FM_F3F4_F5_FromMinus_FT_F3F4),
.number3in3(FM_F3F4_F1_FromPlus_FT_F3F4_number),
.read_add3in3(FM_F3F4_F1_FromPlus_FT_F3F4_read_add),
.read_en3in3(FM_F3F4_F1_FromPlus_FT_F3F4_read_en),
.fullmatch3in3(FM_F3F4_F1_FromPlus_FT_F3F4),
.number4in3(FM_F3F4_F2_FromPlus_FT_F3F4_number),
.read_add4in3(FM_F3F4_F2_FromPlus_FT_F3F4_read_add),
.read_en4in3(FM_F3F4_F2_FromPlus_FT_F3F4_read_en),
.fullmatch4in3(FM_F3F4_F2_FromPlus_FT_F3F4),
.number5in3(FM_F3F4_F5_FromPlus_FT_F3F4_number),
.read_add5in3(FM_F3F4_F5_FromPlus_FT_F3F4_read_add),
.read_en5in3(FM_F3F4_F5_FromPlus_FT_F3F4_read_en),
.fullmatch5in3(FM_F3F4_F5_FromPlus_FT_F3F4),
.trackout(FT_F3F4_TF_F3F4),
.valid_fit(FT_F3F4_TF_F3F4_wr_en),
.start(FM_F3F4_F5_FromPlus_start),
.done(FT_F3F4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

PurgeDuplicate  PD(
.read_add_trackin1(TF_F1F2_PD_read_add),
.trackin1(TF_F1F2_PD),
.read_add_trackin2(TF_F3F4_PD_read_add),
.trackin2(TF_F3F4_PD),
.trackout1(PD_CT_F1F2),
.trackout2(PD_CT_F3F4),
.start(TF_F1F2_start),
.done(PD_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [31:0] reader_out;

wire InputLink_R1Link1_io_rd_ack , InputLink_R1Link2_io_rd_ack , InputLink_R1Link3_io_rd_ack;
wire TPars_L1L2_io_rd_ack , TPars_L3L4_io_rd_ack , TPars_L5L6_io_rd_ack;
// readback mux
// If a particular block is addressed, connect that block's signals
// to the 'rdbk' output. At the same time, assert 'rdbk_sel' to tell downstream muxes to
// use the 'rdbk' from this module as their source of data.
reg [31:0] io_rd_data_reg;
assign io_rd_data = io_rd_data_reg;
// Assert 'io_rd_ack' if any module is asserting its 'rd_ack'.
reg io_rd_ack_reg;
assign io_rd_ack = io_rd_ack_reg;
always @ (posedge io_clk) begin
io_rd_ack_reg <= InputLink_R1Link1_io_rd_ack | InputLink_R1Link2_io_rd_ack | InputLink_R1Link3_io_rd_ack |
TPars_L1L2_io_rd_ack | TPars_L3L4_io_rd_ack | TPars_L5L6_io_rd_ack;
end
// Route the selected register to the 'rdbk' output.
always @(posedge io_clk) begin
if (InputLink_R1Link1_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link1_io_rd_data[31:0];
if (InputLink_R1Link2_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link2_io_rd_data[31:0];
if (InputLink_R1Link3_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link3_io_rd_data[31:0];
if (TPars_L1L2_io_sel) io_rd_data_reg[31:0] <= TPars_L1L2_io_rd_data[31:0];
if (TPars_L3L4_io_sel) io_rd_data_reg[31:0] <= TPars_L3L4_io_rd_data[31:0];
if (TPars_L5L6_io_sel) io_rd_data_reg[31:0] <= TPars_L5L6_io_rd_data[31:0];
//if (reader_ack)    io_rd_data_reg <= reader_out;
end

endmodule
