`timescale 1ns / 1ps

//---------------------------------------------------
// 
//---------------------------------------------------

module spaceinputs(
    
    // inputs
    input clk,
    input reset,
    input BC0,
    input datain,
    input eventin,
    input bxin,
    input numin,
    // outputs
    output dataout
);
    
    always @(posedge clk) begin
        
    end 
      
endmodule
