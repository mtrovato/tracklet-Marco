`timescale 1ns / 1ps
`include "constants.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 09/28/2014 11:01:39 AM
// Design Name:
// Module Name: Tracklet_processing
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module Tracklet_processing(
input clk,
input reset,
input en_proc,
// programming interface
// inputs
input wire io_clk,                    // programming clock
input wire io_sel,                    // this module has been selected for an I/O operation
input wire io_sync,
// start the I/O operation
input wire [15:0] io_addr,        // slave address, memory or register. Top 12 bits already consumed.
input wire io_rd_en,                // this is a read operation
input wire io_wr_en,                // this is a write operation
input wire [31:0] io_wr_data,    // data to write for write operations
// outputs
output wire [31:0] io_rd_data,    // data returned for read operations
output wire io_rd_ack,                // 'read' data from this module is ready
//clocks
input wire [2:0] BX,
input wire first_clk,
input wire not_first_clk,
// inputs
input [31:0] input_link1_reg1,
input [31:0] input_link1_reg2,
input [31:0] input_link2_reg1,
input [31:0] input_link2_reg2,
input [31:0] input_link3_reg1,
input [31:0] input_link3_reg2,
input [31:0] input_link4_reg1,
input [31:0] input_link4_reg2,
input [31:0] input_link5_reg1,
input [31:0] input_link5_reg2,
input [31:0] input_link6_reg1,
input [31:0] input_link6_reg2,
// outputs
input [15:0] BRAM_OUTPUT_addr, // 1 for now, add more later
input BRAM_OUTPUT_clk,
input [31:0] BRAM_OUTPUT_din,
output [31:0] BRAM_OUTPUT_dout,
input BRAM_OUTPUT_en,
input BRAM_OUTPUT_rst,
input [3:0] BRAM_OUTPUT_we,
// Projections L1L2
output wire [50:0] PT_L1L2_Plus_To_DataStream,
output wire PT_L1L2_Plus_To_DataStream_en,
output wire [50:0] PT_L1L2_Minus_To_DataStream,
output wire PT_L1L2_Minus_To_DataStream_en,
input wire [50:0] PT_L1L2_Plus_From_DataStream,
input wire PT_L1L2_Plus_From_DataStream_en,
input wire [50:0] PT_L1L2_Minus_From_DataStream,
input wire PT_L1L2_Minus_From_DataStream_en,
// Projections L3L4
output wire [50:0] PT_L3L4_Plus_To_DataStream,
output wire PT_L3L4_Plus_To_DataStream_en,
output wire [50:0] PT_L3L4_Minus_To_DataStream,
output wire PT_L3L4_Minus_To_DataStream_en,
input wire [50:0] PT_L3L4_Plus_From_DataStream,
input wire PT_L3L4_Plus_From_DataStream_en,
input wire [50:0] PT_L3L4_Minus_From_DataStream,
input wire PT_L3L4_Minus_From_DataStream_en,
// Projections L5L6
output wire [50:0] PT_L5L6_Plus_To_DataStream,
output wire PT_L5L6_Plus_To_DataStream_en,
output wire [50:0] PT_L5L6_Minus_To_DataStream,
output wire PT_L5L6_Minus_To_DataStream_en,
input wire [50:0] PT_L5L6_Plus_From_DataStream,
input wire PT_L5L6_Plus_From_DataStream_en,
input wire [50:0] PT_L5L6_Minus_From_DataStream,
input wire PT_L5L6_Minus_From_DataStream_en,
// Matches L1L2
output wire [38:0] MT_L1L2_Plus_To_DataStream,
output wire MT_L1L2_Plus_To_DataStream_en,
output wire [38:0] MT_L1L2_Minus_To_DataStream,
output wire MT_L1L2_Minus_To_DataStream_en,
input wire [38:0] MT_L1L2_Plus_From_DataStream,
input wire MT_L1L2_Plus_From_DataStream_en,
input wire [38:0] MT_L1L2_Minus_From_DataStream,
input wire MT_L1L2_Minus_From_DataStream_en,
// Matches L3L4
output wire [38:0] MT_L3L4_Plus_To_DataStream,
output wire MT_L3L4_Plus_To_DataStream_en,
output wire [38:0] MT_L3L4_Minus_To_DataStream,
output wire MT_L3L4_Minus_To_DataStream_en,
input wire [38:0] MT_L3L4_Plus_From_DataStream,
input wire MT_L3L4_Plus_From_DataStream_en,
input wire [38:0] MT_L3L4_Minus_From_DataStream,
input wire MT_L3L4_Minus_From_DataStream_en,
// Matches L5L6
output wire [38:0] MT_L5L6_Plus_To_DataStream,
output wire MT_L5L6_Plus_To_DataStream_en,
output wire [38:0] MT_L5L6_Minus_To_DataStream,
output wire MT_L5L6_Minus_To_DataStream_en,
input wire [38:0] MT_L5L6_Plus_From_DataStream,
input wire MT_L5L6_Plus_From_DataStream_en,
input wire [38:0] MT_L5L6_Minus_From_DataStream,
input wire MT_L5L6_Minus_From_DataStream_en,
// Track Fits
output wire [125:0] TF_L1L2_DataStream,
output wire [125:0] TF_L3L4_DataStream,
output wire [125:0] TF_L5L6_DataStream,
output wire [125:0] TF_F1F2_DataStream,
output wire [125:0] TF_F3F4_DataStream

);

// Address bits "io_addr[31:30] = 2'b01" are consumed when selecting 'slave6'
// Address bits "io_addr[29:28] = 2'b01" are consumed when selecting 'tracklet_processing'
wire InputLink_R1Link1_io_sel, TPars_L1L2_io_sel;
wire InputLink_R1Link2_io_sel, TPars_L3L4_io_sel;
wire InputLink_R1Link3_io_sel, TPars_L5L6_io_sel;
wire io_sel_R3_io_block;
assign InputLink_R1Link1_io_sel = io_sel && (io_addr[13:10] == 4'b0001);
assign InputLink_R1Link2_io_sel = io_sel && (io_addr[13:10] == 4'b0010);
assign InputLink_R1Link3_io_sel = io_sel && (io_addr[13:10] == 4'b0011);
assign TPars_L1L2_io_sel  = io_sel && (io_addr[13:10] == 4'b0100);
assign TPars_L3L4_io_sel  = io_sel && (io_addr[13:10] == 4'b0101);
assign TPars_L5L6_io_sel  = io_sel && (io_addr[13:10] == 4'b0110);
assign io_sel_R3_io_block = io_sel && (io_addr[13:10] == 4'b1000);
// data busses for readback
wire [31:0] InputLink_R1Link1_io_rd_data, TPars_L1L2_io_rd_data;
wire [31:0] InputLink_R1Link2_io_rd_data, TPars_L3L4_io_rd_data;
wire [31:0] InputLink_R1Link3_io_rd_data, TPars_L5L6_io_rd_data;

wire IL1_D3_LR1_D3_empty;
wire IL2_D3_LR2_D3_empty;
wire IL3_D3_LR3_D3_empty;

reg [5:0] clk_cnt;

//wire enable_gen;
//enable_generator en_gen(
//.clk(clk),
//.in( (~IL1_D3_LR1_D3_empty | ~IL2_D3_LR2_D3_empty | ~IL3_D3_LR3_D3_empty) & bc0_i ),
//.out(enable_gen)
//);

initial
clk_cnt = 6'b0;
always @(posedge clk) begin
if(en_proc)
clk_cnt <= clk_cnt + 1'b1;
else begin
clk_cnt <= 6'b0;
end
if(clk_cnt == (`tmux - 1'b1))
clk_cnt <= 6'b0;
end

wire [1:0] start1_0, start2_0, start3_0, start4_0, start5_0, startproj5_0, start6_0, start7_0, start8_0, start9_0, start10_0, start11_0;
wire [1:0] done1_0, done2_0, done3_0, done4_0, done_proj4_0, done5_0, done6_0, done7_0, done8_0, done9_0, done10_0;
wire [1:0] start1_5, start2_5, start3_5, start4_5, start5_5, start6_5, start7_5, start8_5, start9_5, start10_5;
wire [1:0] done1_5, done2_5, done3_5, done4_5, done5_5, done6_5, done7_5, done8_5, done9_5, done10_5;

//assign start1_0 = (clk_cnt == 6'd0 && en_proc);
assign start2_0 = done1_0;
assign start3_0 = done2_0;
assign start4_0 = done3_0;
assign start5_0 = done4_0;
assign startproj5_0 = done_proj4_0;
assign start6_0 = done5_0;
assign start7_0 = done6_0;
assign start8_0 = done7_0;
assign start9_0 = done8_0;
assign start10_0 = done9_0;
assign start11_0 = done10_0;

assign start1_5[1] = reset;    // use the top bit of start as reset
assign start1_5[0] = (clk_cnt == 6'd0 && en_proc);
//assign start1_5 = en_proc;
assign start2_5 = done1_5;
assign start3_5 = done2_5;
assign start4_5 = done3_5;
assign start5_5 = done4_5;
assign start6_5 = done5_5;
assign start7_5 = done6_5;
assign start8_5 = done7_5;
assign start9_5 = done8_5;
assign start10_5 = done9_5;




wire IL1_D3_LR1_D3_read_en;
wire [35:0] IL1_D3_LR1_D3;
//wire IL1_D3_LR1_D3_empty;
InputLink  IL1_D3(
.data_in1(input_link1_reg1),
.data_in2(input_link1_reg2),
.read_en(IL1_D3_LR1_D3_read_en),
.data_out(IL1_D3_LR1_D3),
.empty(IL1_D3_LR1_D3_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire IL2_D3_LR2_D3_read_en;
wire [35:0] IL2_D3_LR2_D3;
//wire IL2_D3_LR2_D3_empty;
InputLink  IL2_D3(
.data_in1(input_link2_reg1),
.data_in2(input_link2_reg2),
.read_en(IL2_D3_LR2_D3_read_en),
.data_out(IL2_D3_LR2_D3),
.empty(IL2_D3_LR2_D3_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire IL3_D3_LR3_D3_read_en;
wire [35:0] IL3_D3_LR3_D3;
//wire IL3_D3_LR3_D3_empty;
InputLink  IL3_D3(
.data_in1(input_link3_reg1),
.data_in2(input_link3_reg2),
.read_en(IL3_D3_LR3_D3_read_en),
.data_out(IL3_D3_LR3_D3),
.empty(IL3_D3_LR3_D3_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire IL1_D4_LR1_D4_read_en;
wire [35:0] IL1_D4_LR1_D4;
//wire IL1_D4_LR1_D4_empty;
InputLink  IL1_D4(
.data_in1(input_link4_reg1),
.data_in2(input_link4_reg2),
.read_en(IL1_D4_LR1_D4_read_en),
.data_out(IL1_D4_LR1_D4),
.empty(IL1_D4_LR1_D4_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire IL2_D4_LR2_D4_read_en;
wire [35:0] IL2_D4_LR2_D4;
//wire IL2_D4_LR2_D4_empty;
InputLink  IL2_D4(
.data_in1(input_link5_reg1),
.data_in2(input_link5_reg2),
.read_en(IL2_D4_LR2_D4_read_en),
.data_out(IL2_D4_LR2_D4),
.empty(IL2_D4_LR2_D4_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire IL3_D4_LR3_D4_read_en;
wire [35:0] IL3_D4_LR3_D4;
//wire IL3_D4_LR3_D4_empty;
InputLink  IL3_D4(
.data_in1(input_link6_reg1),
.data_in2(input_link6_reg2),
.read_en(IL3_D4_LR3_D4_read_en),
.data_out(IL3_D4_LR3_D4),
.empty(IL3_D4_LR3_D4_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D3_SL1_L1D3;
wire LR1_D3_SL1_L1D3_wr_en;
wire [5:0] SL1_L1D3_VMR_L1D3_number;
wire [8:0] SL1_L1D3_VMR_L1D3_read_add;
wire [35:0] SL1_L1D3_VMR_L1D3;
StubsByLayer  SL1_L1D3(
.data_in(LR1_D3_SL1_L1D3),
.enable(LR1_D3_SL1_L1D3_wr_en),
.number_out(SL1_L1D3_VMR_L1D3_number),
.read_add(SL1_L1D3_VMR_L1D3_read_add),
.data_out(SL1_L1D3_VMR_L1D3),
.start(start2_0),
.done(done1_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D3_SL2_L1D3;
wire LR2_D3_SL2_L1D3_wr_en;
wire [5:0] SL2_L1D3_VMR_L1D3_number;
wire [8:0] SL2_L1D3_VMR_L1D3_read_add;
wire [35:0] SL2_L1D3_VMR_L1D3;
StubsByLayer  SL2_L1D3(
.data_in(LR2_D3_SL2_L1D3),
.enable(LR2_D3_SL2_L1D3_wr_en),
.number_out(SL2_L1D3_VMR_L1D3_number),
.read_add(SL2_L1D3_VMR_L1D3_read_add),
.data_out(SL2_L1D3_VMR_L1D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D3_SL3_L1D3;
wire LR3_D3_SL3_L1D3_wr_en;
wire [5:0] SL3_L1D3_VMR_L1D3_number;
wire [8:0] SL3_L1D3_VMR_L1D3_read_add;
wire [35:0] SL3_L1D3_VMR_L1D3;
StubsByLayer  SL3_L1D3(
.data_in(LR3_D3_SL3_L1D3),
.enable(LR3_D3_SL3_L1D3_wr_en),
.number_out(SL3_L1D3_VMR_L1D3_number),
.read_add(SL3_L1D3_VMR_L1D3_read_add),
.data_out(SL3_L1D3_VMR_L1D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D4_SL1_L1D4;
wire LR1_D4_SL1_L1D4_wr_en;
wire [5:0] SL1_L1D4_VMR_L1D4_number;
wire [8:0] SL1_L1D4_VMR_L1D4_read_add;
wire [35:0] SL1_L1D4_VMR_L1D4;
StubsByLayer  SL1_L1D4(
.data_in(LR1_D4_SL1_L1D4),
.enable(LR1_D4_SL1_L1D4_wr_en),
.number_out(SL1_L1D4_VMR_L1D4_number),
.read_add(SL1_L1D4_VMR_L1D4_read_add),
.data_out(SL1_L1D4_VMR_L1D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D4_SL2_L1D4;
wire LR2_D4_SL2_L1D4_wr_en;
wire [5:0] SL2_L1D4_VMR_L1D4_number;
wire [8:0] SL2_L1D4_VMR_L1D4_read_add;
wire [35:0] SL2_L1D4_VMR_L1D4;
StubsByLayer  SL2_L1D4(
.data_in(LR2_D4_SL2_L1D4),
.enable(LR2_D4_SL2_L1D4_wr_en),
.number_out(SL2_L1D4_VMR_L1D4_number),
.read_add(SL2_L1D4_VMR_L1D4_read_add),
.data_out(SL2_L1D4_VMR_L1D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D4_SL3_L1D4;
wire LR3_D4_SL3_L1D4_wr_en;
wire [5:0] SL3_L1D4_VMR_L1D4_number;
wire [8:0] SL3_L1D4_VMR_L1D4_read_add;
wire [35:0] SL3_L1D4_VMR_L1D4;
StubsByLayer  SL3_L1D4(
.data_in(LR3_D4_SL3_L1D4),
.enable(LR3_D4_SL3_L1D4_wr_en),
.number_out(SL3_L1D4_VMR_L1D4_number),
.read_add(SL3_L1D4_VMR_L1D4_read_add),
.data_out(SL3_L1D4_VMR_L1D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D3_SL1_L3D3;
wire LR1_D3_SL1_L3D3_wr_en;
wire [5:0] SL1_L3D3_VMR_L3D3_number;
wire [8:0] SL1_L3D3_VMR_L3D3_read_add;
wire [35:0] SL1_L3D3_VMR_L3D3;
StubsByLayer  SL1_L3D3(
.data_in(LR1_D3_SL1_L3D3),
.enable(LR1_D3_SL1_L3D3_wr_en),
.number_out(SL1_L3D3_VMR_L3D3_number),
.read_add(SL1_L3D3_VMR_L3D3_read_add),
.data_out(SL1_L3D3_VMR_L3D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D3_SL2_L3D3;
wire LR2_D3_SL2_L3D3_wr_en;
wire [5:0] SL2_L3D3_VMR_L3D3_number;
wire [8:0] SL2_L3D3_VMR_L3D3_read_add;
wire [35:0] SL2_L3D3_VMR_L3D3;
StubsByLayer  SL2_L3D3(
.data_in(LR2_D3_SL2_L3D3),
.enable(LR2_D3_SL2_L3D3_wr_en),
.number_out(SL2_L3D3_VMR_L3D3_number),
.read_add(SL2_L3D3_VMR_L3D3_read_add),
.data_out(SL2_L3D3_VMR_L3D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D3_SL3_L3D3;
wire LR3_D3_SL3_L3D3_wr_en;
wire [5:0] SL3_L3D3_VMR_L3D3_number;
wire [8:0] SL3_L3D3_VMR_L3D3_read_add;
wire [35:0] SL3_L3D3_VMR_L3D3;
StubsByLayer  SL3_L3D3(
.data_in(LR3_D3_SL3_L3D3),
.enable(LR3_D3_SL3_L3D3_wr_en),
.number_out(SL3_L3D3_VMR_L3D3_number),
.read_add(SL3_L3D3_VMR_L3D3_read_add),
.data_out(SL3_L3D3_VMR_L3D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D4_SL1_L3D4;
wire LR1_D4_SL1_L3D4_wr_en;
wire [5:0] SL1_L3D4_VMR_L3D4_number;
wire [8:0] SL1_L3D4_VMR_L3D4_read_add;
wire [35:0] SL1_L3D4_VMR_L3D4;
StubsByLayer  SL1_L3D4(
.data_in(LR1_D4_SL1_L3D4),
.enable(LR1_D4_SL1_L3D4_wr_en),
.number_out(SL1_L3D4_VMR_L3D4_number),
.read_add(SL1_L3D4_VMR_L3D4_read_add),
.data_out(SL1_L3D4_VMR_L3D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D4_SL2_L3D4;
wire LR2_D4_SL2_L3D4_wr_en;
wire [5:0] SL2_L3D4_VMR_L3D4_number;
wire [8:0] SL2_L3D4_VMR_L3D4_read_add;
wire [35:0] SL2_L3D4_VMR_L3D4;
StubsByLayer  SL2_L3D4(
.data_in(LR2_D4_SL2_L3D4),
.enable(LR2_D4_SL2_L3D4_wr_en),
.number_out(SL2_L3D4_VMR_L3D4_number),
.read_add(SL2_L3D4_VMR_L3D4_read_add),
.data_out(SL2_L3D4_VMR_L3D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D4_SL3_L3D4;
wire LR3_D4_SL3_L3D4_wr_en;
wire [5:0] SL3_L3D4_VMR_L3D4_number;
wire [8:0] SL3_L3D4_VMR_L3D4_read_add;
wire [35:0] SL3_L3D4_VMR_L3D4;
StubsByLayer  SL3_L3D4(
.data_in(LR3_D4_SL3_L3D4),
.enable(LR3_D4_SL3_L3D4_wr_en),
.number_out(SL3_L3D4_VMR_L3D4_number),
.read_add(SL3_L3D4_VMR_L3D4_read_add),
.data_out(SL3_L3D4_VMR_L3D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D3_SL1_L5D3;
wire LR1_D3_SL1_L5D3_wr_en;
wire [5:0] SL1_L5D3_VMR_L5D3_number;
wire [8:0] SL1_L5D3_VMR_L5D3_read_add;
wire [35:0] SL1_L5D3_VMR_L5D3;
StubsByLayer  SL1_L5D3(
.data_in(LR1_D3_SL1_L5D3),
.enable(LR1_D3_SL1_L5D3_wr_en),
.number_out(SL1_L5D3_VMR_L5D3_number),
.read_add(SL1_L5D3_VMR_L5D3_read_add),
.data_out(SL1_L5D3_VMR_L5D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D3_SL2_L5D3;
wire LR2_D3_SL2_L5D3_wr_en;
wire [5:0] SL2_L5D3_VMR_L5D3_number;
wire [8:0] SL2_L5D3_VMR_L5D3_read_add;
wire [35:0] SL2_L5D3_VMR_L5D3;
StubsByLayer  SL2_L5D3(
.data_in(LR2_D3_SL2_L5D3),
.enable(LR2_D3_SL2_L5D3_wr_en),
.number_out(SL2_L5D3_VMR_L5D3_number),
.read_add(SL2_L5D3_VMR_L5D3_read_add),
.data_out(SL2_L5D3_VMR_L5D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D3_SL3_L5D3;
wire LR3_D3_SL3_L5D3_wr_en;
wire [5:0] SL3_L5D3_VMR_L5D3_number;
wire [8:0] SL3_L5D3_VMR_L5D3_read_add;
wire [35:0] SL3_L5D3_VMR_L5D3;
StubsByLayer  SL3_L5D3(
.data_in(LR3_D3_SL3_L5D3),
.enable(LR3_D3_SL3_L5D3_wr_en),
.number_out(SL3_L5D3_VMR_L5D3_number),
.read_add(SL3_L5D3_VMR_L5D3_read_add),
.data_out(SL3_L5D3_VMR_L5D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D4_SL1_L5D4;
wire LR1_D4_SL1_L5D4_wr_en;
wire [5:0] SL1_L5D4_VMR_L5D4_number;
wire [8:0] SL1_L5D4_VMR_L5D4_read_add;
wire [35:0] SL1_L5D4_VMR_L5D4;
StubsByLayer  SL1_L5D4(
.data_in(LR1_D4_SL1_L5D4),
.enable(LR1_D4_SL1_L5D4_wr_en),
.number_out(SL1_L5D4_VMR_L5D4_number),
.read_add(SL1_L5D4_VMR_L5D4_read_add),
.data_out(SL1_L5D4_VMR_L5D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D4_SL2_L5D4;
wire LR2_D4_SL2_L5D4_wr_en;
wire [5:0] SL2_L5D4_VMR_L5D4_number;
wire [8:0] SL2_L5D4_VMR_L5D4_read_add;
wire [35:0] SL2_L5D4_VMR_L5D4;
StubsByLayer  SL2_L5D4(
.data_in(LR2_D4_SL2_L5D4),
.enable(LR2_D4_SL2_L5D4_wr_en),
.number_out(SL2_L5D4_VMR_L5D4_number),
.read_add(SL2_L5D4_VMR_L5D4_read_add),
.data_out(SL2_L5D4_VMR_L5D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D4_SL3_L5D4;
wire LR3_D4_SL3_L5D4_wr_en;
wire [5:0] SL3_L5D4_VMR_L5D4_number;
wire [8:0] SL3_L5D4_VMR_L5D4_read_add;
wire [35:0] SL3_L5D4_VMR_L5D4;
StubsByLayer  SL3_L5D4(
.data_in(LR3_D4_SL3_L5D4),
.enable(LR3_D4_SL3_L5D4_wr_en),
.number_out(SL3_L5D4_VMR_L5D4_number),
.read_add(SL3_L5D4_VMR_L5D4_read_add),
.data_out(SL3_L5D4_VMR_L5D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D3_SL1_L2D3;
wire LR1_D3_SL1_L2D3_wr_en;
wire [5:0] SL1_L2D3_VMR_L2D3_number;
wire [8:0] SL1_L2D3_VMR_L2D3_read_add;
wire [35:0] SL1_L2D3_VMR_L2D3;
StubsByLayer  SL1_L2D3(
.data_in(LR1_D3_SL1_L2D3),
.enable(LR1_D3_SL1_L2D3_wr_en),
.number_out(SL1_L2D3_VMR_L2D3_number),
.read_add(SL1_L2D3_VMR_L2D3_read_add),
.data_out(SL1_L2D3_VMR_L2D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D3_SL2_L2D3;
wire LR2_D3_SL2_L2D3_wr_en;
wire [5:0] SL2_L2D3_VMR_L2D3_number;
wire [8:0] SL2_L2D3_VMR_L2D3_read_add;
wire [35:0] SL2_L2D3_VMR_L2D3;
StubsByLayer  SL2_L2D3(
.data_in(LR2_D3_SL2_L2D3),
.enable(LR2_D3_SL2_L2D3_wr_en),
.number_out(SL2_L2D3_VMR_L2D3_number),
.read_add(SL2_L2D3_VMR_L2D3_read_add),
.data_out(SL2_L2D3_VMR_L2D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D3_SL3_L2D3;
wire LR3_D3_SL3_L2D3_wr_en;
wire [5:0] SL3_L2D3_VMR_L2D3_number;
wire [8:0] SL3_L2D3_VMR_L2D3_read_add;
wire [35:0] SL3_L2D3_VMR_L2D3;
StubsByLayer  SL3_L2D3(
.data_in(LR3_D3_SL3_L2D3),
.enable(LR3_D3_SL3_L2D3_wr_en),
.number_out(SL3_L2D3_VMR_L2D3_number),
.read_add(SL3_L2D3_VMR_L2D3_read_add),
.data_out(SL3_L2D3_VMR_L2D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D4_SL1_L2D4;
wire LR1_D4_SL1_L2D4_wr_en;
wire [5:0] SL1_L2D4_VMR_L2D4_number;
wire [8:0] SL1_L2D4_VMR_L2D4_read_add;
wire [35:0] SL1_L2D4_VMR_L2D4;
StubsByLayer  SL1_L2D4(
.data_in(LR1_D4_SL1_L2D4),
.enable(LR1_D4_SL1_L2D4_wr_en),
.number_out(SL1_L2D4_VMR_L2D4_number),
.read_add(SL1_L2D4_VMR_L2D4_read_add),
.data_out(SL1_L2D4_VMR_L2D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D4_SL2_L2D4;
wire LR2_D4_SL2_L2D4_wr_en;
wire [5:0] SL2_L2D4_VMR_L2D4_number;
wire [8:0] SL2_L2D4_VMR_L2D4_read_add;
wire [35:0] SL2_L2D4_VMR_L2D4;
StubsByLayer  SL2_L2D4(
.data_in(LR2_D4_SL2_L2D4),
.enable(LR2_D4_SL2_L2D4_wr_en),
.number_out(SL2_L2D4_VMR_L2D4_number),
.read_add(SL2_L2D4_VMR_L2D4_read_add),
.data_out(SL2_L2D4_VMR_L2D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D4_SL3_L2D4;
wire LR3_D4_SL3_L2D4_wr_en;
wire [5:0] SL3_L2D4_VMR_L2D4_number;
wire [8:0] SL3_L2D4_VMR_L2D4_read_add;
wire [35:0] SL3_L2D4_VMR_L2D4;
StubsByLayer  SL3_L2D4(
.data_in(LR3_D4_SL3_L2D4),
.enable(LR3_D4_SL3_L2D4_wr_en),
.number_out(SL3_L2D4_VMR_L2D4_number),
.read_add(SL3_L2D4_VMR_L2D4_read_add),
.data_out(SL3_L2D4_VMR_L2D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D3_SL1_L4D3;
wire LR1_D3_SL1_L4D3_wr_en;
wire [5:0] SL1_L4D3_VMR_L4D3_number;
wire [8:0] SL1_L4D3_VMR_L4D3_read_add;
wire [35:0] SL1_L4D3_VMR_L4D3;
StubsByLayer  SL1_L4D3(
.data_in(LR1_D3_SL1_L4D3),
.enable(LR1_D3_SL1_L4D3_wr_en),
.number_out(SL1_L4D3_VMR_L4D3_number),
.read_add(SL1_L4D3_VMR_L4D3_read_add),
.data_out(SL1_L4D3_VMR_L4D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D3_SL2_L4D3;
wire LR2_D3_SL2_L4D3_wr_en;
wire [5:0] SL2_L4D3_VMR_L4D3_number;
wire [8:0] SL2_L4D3_VMR_L4D3_read_add;
wire [35:0] SL2_L4D3_VMR_L4D3;
StubsByLayer  SL2_L4D3(
.data_in(LR2_D3_SL2_L4D3),
.enable(LR2_D3_SL2_L4D3_wr_en),
.number_out(SL2_L4D3_VMR_L4D3_number),
.read_add(SL2_L4D3_VMR_L4D3_read_add),
.data_out(SL2_L4D3_VMR_L4D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D3_SL3_L4D3;
wire LR3_D3_SL3_L4D3_wr_en;
wire [5:0] SL3_L4D3_VMR_L4D3_number;
wire [8:0] SL3_L4D3_VMR_L4D3_read_add;
wire [35:0] SL3_L4D3_VMR_L4D3;
StubsByLayer  SL3_L4D3(
.data_in(LR3_D3_SL3_L4D3),
.enable(LR3_D3_SL3_L4D3_wr_en),
.number_out(SL3_L4D3_VMR_L4D3_number),
.read_add(SL3_L4D3_VMR_L4D3_read_add),
.data_out(SL3_L4D3_VMR_L4D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D4_SL1_L4D4;
wire LR1_D4_SL1_L4D4_wr_en;
wire [5:0] SL1_L4D4_VMR_L4D4_number;
wire [8:0] SL1_L4D4_VMR_L4D4_read_add;
wire [35:0] SL1_L4D4_VMR_L4D4;
StubsByLayer  SL1_L4D4(
.data_in(LR1_D4_SL1_L4D4),
.enable(LR1_D4_SL1_L4D4_wr_en),
.number_out(SL1_L4D4_VMR_L4D4_number),
.read_add(SL1_L4D4_VMR_L4D4_read_add),
.data_out(SL1_L4D4_VMR_L4D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D4_SL2_L4D4;
wire LR2_D4_SL2_L4D4_wr_en;
wire [5:0] SL2_L4D4_VMR_L4D4_number;
wire [8:0] SL2_L4D4_VMR_L4D4_read_add;
wire [35:0] SL2_L4D4_VMR_L4D4;
StubsByLayer  SL2_L4D4(
.data_in(LR2_D4_SL2_L4D4),
.enable(LR2_D4_SL2_L4D4_wr_en),
.number_out(SL2_L4D4_VMR_L4D4_number),
.read_add(SL2_L4D4_VMR_L4D4_read_add),
.data_out(SL2_L4D4_VMR_L4D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D4_SL3_L4D4;
wire LR3_D4_SL3_L4D4_wr_en;
wire [5:0] SL3_L4D4_VMR_L4D4_number;
wire [8:0] SL3_L4D4_VMR_L4D4_read_add;
wire [35:0] SL3_L4D4_VMR_L4D4;
StubsByLayer  SL3_L4D4(
.data_in(LR3_D4_SL3_L4D4),
.enable(LR3_D4_SL3_L4D4_wr_en),
.number_out(SL3_L4D4_VMR_L4D4_number),
.read_add(SL3_L4D4_VMR_L4D4_read_add),
.data_out(SL3_L4D4_VMR_L4D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D3_SL1_L6D3;
wire LR1_D3_SL1_L6D3_wr_en;
wire [5:0] SL1_L6D3_VMR_L6D3_number;
wire [8:0] SL1_L6D3_VMR_L6D3_read_add;
wire [35:0] SL1_L6D3_VMR_L6D3;
StubsByLayer  SL1_L6D3(
.data_in(LR1_D3_SL1_L6D3),
.enable(LR1_D3_SL1_L6D3_wr_en),
.number_out(SL1_L6D3_VMR_L6D3_number),
.read_add(SL1_L6D3_VMR_L6D3_read_add),
.data_out(SL1_L6D3_VMR_L6D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D3_SL2_L6D3;
wire LR2_D3_SL2_L6D3_wr_en;
wire [5:0] SL2_L6D3_VMR_L6D3_number;
wire [8:0] SL2_L6D3_VMR_L6D3_read_add;
wire [35:0] SL2_L6D3_VMR_L6D3;
StubsByLayer  SL2_L6D3(
.data_in(LR2_D3_SL2_L6D3),
.enable(LR2_D3_SL2_L6D3_wr_en),
.number_out(SL2_L6D3_VMR_L6D3_number),
.read_add(SL2_L6D3_VMR_L6D3_read_add),
.data_out(SL2_L6D3_VMR_L6D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D3_SL3_L6D3;
wire LR3_D3_SL3_L6D3_wr_en;
wire [5:0] SL3_L6D3_VMR_L6D3_number;
wire [8:0] SL3_L6D3_VMR_L6D3_read_add;
wire [35:0] SL3_L6D3_VMR_L6D3;
StubsByLayer  SL3_L6D3(
.data_in(LR3_D3_SL3_L6D3),
.enable(LR3_D3_SL3_L6D3_wr_en),
.number_out(SL3_L6D3_VMR_L6D3_number),
.read_add(SL3_L6D3_VMR_L6D3_read_add),
.data_out(SL3_L6D3_VMR_L6D3),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR1_D4_SL1_L6D4;
wire LR1_D4_SL1_L6D4_wr_en;
wire [5:0] SL1_L6D4_VMR_L6D4_number;
wire [8:0] SL1_L6D4_VMR_L6D4_read_add;
wire [35:0] SL1_L6D4_VMR_L6D4;
StubsByLayer  SL1_L6D4(
.data_in(LR1_D4_SL1_L6D4),
.enable(LR1_D4_SL1_L6D4_wr_en),
.number_out(SL1_L6D4_VMR_L6D4_number),
.read_add(SL1_L6D4_VMR_L6D4_read_add),
.data_out(SL1_L6D4_VMR_L6D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR2_D4_SL2_L6D4;
wire LR2_D4_SL2_L6D4_wr_en;
wire [5:0] SL2_L6D4_VMR_L6D4_number;
wire [8:0] SL2_L6D4_VMR_L6D4_read_add;
wire [35:0] SL2_L6D4_VMR_L6D4;
StubsByLayer  SL2_L6D4(
.data_in(LR2_D4_SL2_L6D4),
.enable(LR2_D4_SL2_L6D4_wr_en),
.number_out(SL2_L6D4_VMR_L6D4_number),
.read_add(SL2_L6D4_VMR_L6D4_read_add),
.data_out(SL2_L6D4_VMR_L6D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] LR3_D4_SL3_L6D4;
wire LR3_D4_SL3_L6D4_wr_en;
wire [5:0] SL3_L6D4_VMR_L6D4_number;
wire [8:0] SL3_L6D4_VMR_L6D4_read_add;
wire [35:0] SL3_L6D4_VMR_L6D4;
StubsByLayer  SL3_L6D4(
.data_in(LR3_D4_SL3_L6D4),
.enable(LR3_D4_SL3_L6D4_wr_en),
.number_out(SL3_L6D4_VMR_L6D4_number),
.read_add(SL3_L6D4_VMR_L6D4_read_add),
.data_out(SL3_L6D4_VMR_L6D4),
.start(start2_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z1n1;
wire VMR_L1D3_VMS_L1D3PHI1Z1n1_wr_en;
wire [5:0] VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_number;
wire [10:0] VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_read_add;
wire [17:0] VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1;
VMStubs #("Tracklet") VMS_L1D3PHI1Z1n1(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z1n1),
.enable(VMR_L1D3_VMS_L1D3PHI1Z1n1_wr_en),
.number_out(VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_number),
.read_add(VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_read_add),
.data_out(VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1),
.start(start3_0),
.done(done2_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI1Z1n1;
wire VMR_L2D3_VMS_L2D3PHI1Z1n1_wr_en;
wire [5:0] VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_number;
wire [10:0] VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_read_add;
wire [17:0] VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1;
VMStubs #("Tracklet") VMS_L2D3PHI1Z1n1(
.data_in(VMR_L2D3_VMS_L2D3PHI1Z1n1),
.enable(VMR_L2D3_VMS_L2D3PHI1Z1n1_wr_en),
.number_out(VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_number),
.read_add(VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_read_add),
.data_out(VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z1n2;
wire VMR_L1D3_VMS_L1D3PHI1Z1n2_wr_en;
wire [5:0] VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1_number;
wire [10:0] VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1_read_add;
wire [17:0] VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1;
VMStubs #("Tracklet") VMS_L1D3PHI1Z1n2(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z1n2),
.enable(VMR_L1D3_VMS_L1D3PHI1Z1n2_wr_en),
.number_out(VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1_number),
.read_add(VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1_read_add),
.data_out(VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z1n1;
wire VMR_L2D3_VMS_L2D3PHI2Z1n1_wr_en;
wire [5:0] VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1_number;
wire [10:0] VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1_read_add;
wire [17:0] VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1;
VMStubs #("Tracklet") VMS_L2D3PHI2Z1n1(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z1n1),
.enable(VMR_L2D3_VMS_L2D3PHI2Z1n1_wr_en),
.number_out(VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1_number),
.read_add(VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1_read_add),
.data_out(VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z1n1;
wire VMR_L1D3_VMS_L1D3PHI2Z1n1_wr_en;
wire [5:0] VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1_number;
wire [10:0] VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1_read_add;
wire [17:0] VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1;
VMStubs #("Tracklet") VMS_L1D3PHI2Z1n1(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z1n1),
.enable(VMR_L1D3_VMS_L1D3PHI2Z1n1_wr_en),
.number_out(VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1_number),
.read_add(VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1_read_add),
.data_out(VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z1n2;
wire VMR_L2D3_VMS_L2D3PHI2Z1n2_wr_en;
wire [5:0] VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1_number;
wire [10:0] VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1_read_add;
wire [17:0] VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1;
VMStubs #("Tracklet") VMS_L2D3PHI2Z1n2(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z1n2),
.enable(VMR_L2D3_VMS_L2D3PHI2Z1n2_wr_en),
.number_out(VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1_number),
.read_add(VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1_read_add),
.data_out(VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z1n2;
wire VMR_L1D3_VMS_L1D3PHI2Z1n2_wr_en;
wire [5:0] VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1_number;
wire [10:0] VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1_read_add;
wire [17:0] VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1;
VMStubs #("Tracklet") VMS_L1D3PHI2Z1n2(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z1n2),
.enable(VMR_L1D3_VMS_L1D3PHI2Z1n2_wr_en),
.number_out(VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1_number),
.read_add(VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1_read_add),
.data_out(VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z1n1;
wire VMR_L2D3_VMS_L2D3PHI3Z1n1_wr_en;
wire [5:0] VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1_number;
wire [10:0] VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1_read_add;
wire [17:0] VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1;
VMStubs #("Tracklet") VMS_L2D3PHI3Z1n1(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z1n1),
.enable(VMR_L2D3_VMS_L2D3PHI3Z1n1_wr_en),
.number_out(VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1_number),
.read_add(VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1_read_add),
.data_out(VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z1n1;
wire VMR_L1D3_VMS_L1D3PHI3Z1n1_wr_en;
wire [5:0] VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1_number;
wire [10:0] VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1_read_add;
wire [17:0] VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1;
VMStubs #("Tracklet") VMS_L1D3PHI3Z1n1(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z1n1),
.enable(VMR_L1D3_VMS_L1D3PHI3Z1n1_wr_en),
.number_out(VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1_number),
.read_add(VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1_read_add),
.data_out(VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z1n2;
wire VMR_L2D3_VMS_L2D3PHI3Z1n2_wr_en;
wire [5:0] VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1_number;
wire [10:0] VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1_read_add;
wire [17:0] VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1;
VMStubs #("Tracklet") VMS_L2D3PHI3Z1n2(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z1n2),
.enable(VMR_L2D3_VMS_L2D3PHI3Z1n2_wr_en),
.number_out(VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1_number),
.read_add(VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1_read_add),
.data_out(VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z1n2;
wire VMR_L1D3_VMS_L1D3PHI3Z1n2_wr_en;
wire [5:0] VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1_number;
wire [10:0] VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1_read_add;
wire [17:0] VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1;
VMStubs #("Tracklet") VMS_L1D3PHI3Z1n2(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z1n2),
.enable(VMR_L1D3_VMS_L1D3PHI3Z1n2_wr_en),
.number_out(VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1_number),
.read_add(VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1_read_add),
.data_out(VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI4Z1n1;
wire VMR_L2D3_VMS_L2D3PHI4Z1n1_wr_en;
wire [5:0] VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1_number;
wire [10:0] VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1_read_add;
wire [17:0] VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1;
VMStubs #("Tracklet") VMS_L2D3PHI4Z1n1(
.data_in(VMR_L2D3_VMS_L2D3PHI4Z1n1),
.enable(VMR_L2D3_VMS_L2D3PHI4Z1n1_wr_en),
.number_out(VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1_number),
.read_add(VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1_read_add),
.data_out(VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z1n3;
wire VMR_L1D3_VMS_L1D3PHI1Z1n3_wr_en;
wire [5:0] VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2_number;
wire [10:0] VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2_read_add;
wire [17:0] VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2;
VMStubs #("Tracklet") VMS_L1D3PHI1Z1n3(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z1n3),
.enable(VMR_L1D3_VMS_L1D3PHI1Z1n3_wr_en),
.number_out(VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2_number),
.read_add(VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2_read_add),
.data_out(VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI1Z2n1;
wire VMR_L2D3_VMS_L2D3PHI1Z2n1_wr_en;
wire [5:0] VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2_number;
wire [10:0] VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2_read_add;
wire [17:0] VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2;
VMStubs #("Tracklet") VMS_L2D3PHI1Z2n1(
.data_in(VMR_L2D3_VMS_L2D3PHI1Z2n1),
.enable(VMR_L2D3_VMS_L2D3PHI1Z2n1_wr_en),
.number_out(VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2_number),
.read_add(VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2_read_add),
.data_out(VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z1n4;
wire VMR_L1D3_VMS_L1D3PHI1Z1n4_wr_en;
wire [5:0] VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2_number;
wire [10:0] VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2;
VMStubs #("Tracklet") VMS_L1D3PHI1Z1n4(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z1n4),
.enable(VMR_L1D3_VMS_L1D3PHI1Z1n4_wr_en),
.number_out(VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2_number),
.read_add(VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2_read_add),
.data_out(VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z2n1;
wire VMR_L2D3_VMS_L2D3PHI2Z2n1_wr_en;
wire [5:0] VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2_number;
wire [10:0] VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2;
VMStubs #("Tracklet") VMS_L2D3PHI2Z2n1(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z2n1),
.enable(VMR_L2D3_VMS_L2D3PHI2Z2n1_wr_en),
.number_out(VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2_number),
.read_add(VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2_read_add),
.data_out(VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z1n3;
wire VMR_L1D3_VMS_L1D3PHI2Z1n3_wr_en;
wire [5:0] VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2_number;
wire [10:0] VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2;
VMStubs #("Tracklet") VMS_L1D3PHI2Z1n3(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z1n3),
.enable(VMR_L1D3_VMS_L1D3PHI2Z1n3_wr_en),
.number_out(VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2_number),
.read_add(VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2_read_add),
.data_out(VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z2n2;
wire VMR_L2D3_VMS_L2D3PHI2Z2n2_wr_en;
wire [5:0] VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2_number;
wire [10:0] VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2;
VMStubs #("Tracklet") VMS_L2D3PHI2Z2n2(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z2n2),
.enable(VMR_L2D3_VMS_L2D3PHI2Z2n2_wr_en),
.number_out(VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2_number),
.read_add(VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2_read_add),
.data_out(VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z1n4;
wire VMR_L1D3_VMS_L1D3PHI2Z1n4_wr_en;
wire [5:0] VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2_number;
wire [10:0] VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2;
VMStubs #("Tracklet") VMS_L1D3PHI2Z1n4(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z1n4),
.enable(VMR_L1D3_VMS_L1D3PHI2Z1n4_wr_en),
.number_out(VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2_number),
.read_add(VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2_read_add),
.data_out(VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z2n1;
wire VMR_L2D3_VMS_L2D3PHI3Z2n1_wr_en;
wire [5:0] VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2_number;
wire [10:0] VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2;
VMStubs #("Tracklet") VMS_L2D3PHI3Z2n1(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z2n1),
.enable(VMR_L2D3_VMS_L2D3PHI3Z2n1_wr_en),
.number_out(VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2_number),
.read_add(VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2_read_add),
.data_out(VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z1n3;
wire VMR_L1D3_VMS_L1D3PHI3Z1n3_wr_en;
wire [5:0] VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2_number;
wire [10:0] VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2;
VMStubs #("Tracklet") VMS_L1D3PHI3Z1n3(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z1n3),
.enable(VMR_L1D3_VMS_L1D3PHI3Z1n3_wr_en),
.number_out(VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2_number),
.read_add(VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2_read_add),
.data_out(VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z2n2;
wire VMR_L2D3_VMS_L2D3PHI3Z2n2_wr_en;
wire [5:0] VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2_number;
wire [10:0] VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2;
VMStubs #("Tracklet") VMS_L2D3PHI3Z2n2(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z2n2),
.enable(VMR_L2D3_VMS_L2D3PHI3Z2n2_wr_en),
.number_out(VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2_number),
.read_add(VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2_read_add),
.data_out(VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z1n4;
wire VMR_L1D3_VMS_L1D3PHI3Z1n4_wr_en;
wire [5:0] VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2_number;
wire [10:0] VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2_read_add;
wire [17:0] VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2;
VMStubs #("Tracklet") VMS_L1D3PHI3Z1n4(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z1n4),
.enable(VMR_L1D3_VMS_L1D3PHI3Z1n4_wr_en),
.number_out(VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2_number),
.read_add(VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2_read_add),
.data_out(VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI4Z2n1;
wire VMR_L2D3_VMS_L2D3PHI4Z2n1_wr_en;
wire [5:0] VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2_number;
wire [10:0] VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2_read_add;
wire [17:0] VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2;
VMStubs #("Tracklet") VMS_L2D3PHI4Z2n1(
.data_in(VMR_L2D3_VMS_L2D3PHI4Z2n1),
.enable(VMR_L2D3_VMS_L2D3PHI4Z2n1_wr_en),
.number_out(VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2_number),
.read_add(VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2_read_add),
.data_out(VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z2n1;
wire VMR_L1D3_VMS_L1D3PHI1Z2n1_wr_en;
wire [5:0] VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2_number;
wire [10:0] VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2_read_add;
wire [17:0] VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2;
VMStubs #("Tracklet") VMS_L1D3PHI1Z2n1(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z2n1),
.enable(VMR_L1D3_VMS_L1D3PHI1Z2n1_wr_en),
.number_out(VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2_number),
.read_add(VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2_read_add),
.data_out(VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI1Z2n2;
wire VMR_L2D3_VMS_L2D3PHI1Z2n2_wr_en;
wire [5:0] VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2_number;
wire [10:0] VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2_read_add;
wire [17:0] VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2;
VMStubs #("Tracklet") VMS_L2D3PHI1Z2n2(
.data_in(VMR_L2D3_VMS_L2D3PHI1Z2n2),
.enable(VMR_L2D3_VMS_L2D3PHI1Z2n2_wr_en),
.number_out(VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2_number),
.read_add(VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2_read_add),
.data_out(VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z2n2;
wire VMR_L1D3_VMS_L1D3PHI1Z2n2_wr_en;
wire [5:0] VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2_number;
wire [10:0] VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2;
VMStubs #("Tracklet") VMS_L1D3PHI1Z2n2(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z2n2),
.enable(VMR_L1D3_VMS_L1D3PHI1Z2n2_wr_en),
.number_out(VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2_number),
.read_add(VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2_read_add),
.data_out(VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z2n3;
wire VMR_L2D3_VMS_L2D3PHI2Z2n3_wr_en;
wire [5:0] VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2_number;
wire [10:0] VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2;
VMStubs #("Tracklet") VMS_L2D3PHI2Z2n3(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z2n3),
.enable(VMR_L2D3_VMS_L2D3PHI2Z2n3_wr_en),
.number_out(VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2_number),
.read_add(VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2_read_add),
.data_out(VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z2n1;
wire VMR_L1D3_VMS_L1D3PHI2Z2n1_wr_en;
wire [5:0] VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2_number;
wire [10:0] VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2;
VMStubs #("Tracklet") VMS_L1D3PHI2Z2n1(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z2n1),
.enable(VMR_L1D3_VMS_L1D3PHI2Z2n1_wr_en),
.number_out(VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2_number),
.read_add(VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2_read_add),
.data_out(VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z2n4;
wire VMR_L2D3_VMS_L2D3PHI2Z2n4_wr_en;
wire [5:0] VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2_number;
wire [10:0] VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2;
VMStubs #("Tracklet") VMS_L2D3PHI2Z2n4(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z2n4),
.enable(VMR_L2D3_VMS_L2D3PHI2Z2n4_wr_en),
.number_out(VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2_number),
.read_add(VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2_read_add),
.data_out(VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z2n2;
wire VMR_L1D3_VMS_L1D3PHI2Z2n2_wr_en;
wire [5:0] VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2_number;
wire [10:0] VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2;
VMStubs #("Tracklet") VMS_L1D3PHI2Z2n2(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z2n2),
.enable(VMR_L1D3_VMS_L1D3PHI2Z2n2_wr_en),
.number_out(VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2_number),
.read_add(VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2_read_add),
.data_out(VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z2n3;
wire VMR_L2D3_VMS_L2D3PHI3Z2n3_wr_en;
wire [5:0] VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2_number;
wire [10:0] VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2;
VMStubs #("Tracklet") VMS_L2D3PHI3Z2n3(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z2n3),
.enable(VMR_L2D3_VMS_L2D3PHI3Z2n3_wr_en),
.number_out(VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2_number),
.read_add(VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2_read_add),
.data_out(VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z2n1;
wire VMR_L1D3_VMS_L1D3PHI3Z2n1_wr_en;
wire [5:0] VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2_number;
wire [10:0] VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2;
VMStubs #("Tracklet") VMS_L1D3PHI3Z2n1(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z2n1),
.enable(VMR_L1D3_VMS_L1D3PHI3Z2n1_wr_en),
.number_out(VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2_number),
.read_add(VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2_read_add),
.data_out(VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z2n4;
wire VMR_L2D3_VMS_L2D3PHI3Z2n4_wr_en;
wire [5:0] VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2_number;
wire [10:0] VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2;
VMStubs #("Tracklet") VMS_L2D3PHI3Z2n4(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z2n4),
.enable(VMR_L2D3_VMS_L2D3PHI3Z2n4_wr_en),
.number_out(VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2_number),
.read_add(VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2_read_add),
.data_out(VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z2n2;
wire VMR_L1D3_VMS_L1D3PHI3Z2n2_wr_en;
wire [5:0] VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_number;
wire [10:0] VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_read_add;
wire [17:0] VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2;
VMStubs #("Tracklet") VMS_L1D3PHI3Z2n2(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z2n2),
.enable(VMR_L1D3_VMS_L1D3PHI3Z2n2_wr_en),
.number_out(VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_number),
.read_add(VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_read_add),
.data_out(VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI4Z2n2;
wire VMR_L2D3_VMS_L2D3PHI4Z2n2_wr_en;
wire [5:0] VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_number;
wire [10:0] VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_read_add;
wire [17:0] VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2;
VMStubs #("Tracklet") VMS_L2D3PHI4Z2n2(
.data_in(VMR_L2D3_VMS_L2D3PHI4Z2n2),
.enable(VMR_L2D3_VMS_L2D3PHI4Z2n2_wr_en),
.number_out(VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_number),
.read_add(VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_read_add),
.data_out(VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z1n5;
wire VMR_L1D3_VMS_L1D3PHI1Z1n5_wr_en;
wire [5:0] VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1_number;
wire [10:0] VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1_read_add;
wire [17:0] VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1;
VMStubs #("Tracklet") VMS_L1D3PHI1Z1n5(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z1n5),
.enable(VMR_L1D3_VMS_L1D3PHI1Z1n5_wr_en),
.number_out(VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1_number),
.read_add(VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1_read_add),
.data_out(VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI1Z1n1;
wire VMR_L2D4_VMS_L2D4PHI1Z1n1_wr_en;
wire [5:0] VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1_number;
wire [10:0] VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1_read_add;
wire [17:0] VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1;
VMStubs #("Tracklet") VMS_L2D4PHI1Z1n1(
.data_in(VMR_L2D4_VMS_L2D4PHI1Z1n1),
.enable(VMR_L2D4_VMS_L2D4PHI1Z1n1_wr_en),
.number_out(VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1_number),
.read_add(VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1_read_add),
.data_out(VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z1n6;
wire VMR_L1D3_VMS_L1D3PHI1Z1n6_wr_en;
wire [5:0] VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1_number;
wire [10:0] VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1;
VMStubs #("Tracklet") VMS_L1D3PHI1Z1n6(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z1n6),
.enable(VMR_L1D3_VMS_L1D3PHI1Z1n6_wr_en),
.number_out(VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1_number),
.read_add(VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1_read_add),
.data_out(VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z1n1;
wire VMR_L2D4_VMS_L2D4PHI2Z1n1_wr_en;
wire [5:0] VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1_number;
wire [10:0] VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1;
VMStubs #("Tracklet") VMS_L2D4PHI2Z1n1(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z1n1),
.enable(VMR_L2D4_VMS_L2D4PHI2Z1n1_wr_en),
.number_out(VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1_number),
.read_add(VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1_read_add),
.data_out(VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z1n5;
wire VMR_L1D3_VMS_L1D3PHI2Z1n5_wr_en;
wire [5:0] VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1_number;
wire [10:0] VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1;
VMStubs #("Tracklet") VMS_L1D3PHI2Z1n5(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z1n5),
.enable(VMR_L1D3_VMS_L1D3PHI2Z1n5_wr_en),
.number_out(VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1_number),
.read_add(VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1_read_add),
.data_out(VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z1n2;
wire VMR_L2D4_VMS_L2D4PHI2Z1n2_wr_en;
wire [5:0] VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1_number;
wire [10:0] VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1;
VMStubs #("Tracklet") VMS_L2D4PHI2Z1n2(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z1n2),
.enable(VMR_L2D4_VMS_L2D4PHI2Z1n2_wr_en),
.number_out(VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1_number),
.read_add(VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1_read_add),
.data_out(VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z1n6;
wire VMR_L1D3_VMS_L1D3PHI2Z1n6_wr_en;
wire [5:0] VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1_number;
wire [10:0] VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1;
VMStubs #("Tracklet") VMS_L1D3PHI2Z1n6(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z1n6),
.enable(VMR_L1D3_VMS_L1D3PHI2Z1n6_wr_en),
.number_out(VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1_number),
.read_add(VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1_read_add),
.data_out(VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z1n1;
wire VMR_L2D4_VMS_L2D4PHI3Z1n1_wr_en;
wire [5:0] VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1_number;
wire [10:0] VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1;
VMStubs #("Tracklet") VMS_L2D4PHI3Z1n1(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z1n1),
.enable(VMR_L2D4_VMS_L2D4PHI3Z1n1_wr_en),
.number_out(VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1_number),
.read_add(VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1_read_add),
.data_out(VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z1n5;
wire VMR_L1D3_VMS_L1D3PHI3Z1n5_wr_en;
wire [5:0] VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1_number;
wire [10:0] VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1;
VMStubs #("Tracklet") VMS_L1D3PHI3Z1n5(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z1n5),
.enable(VMR_L1D3_VMS_L1D3PHI3Z1n5_wr_en),
.number_out(VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1_number),
.read_add(VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1_read_add),
.data_out(VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z1n2;
wire VMR_L2D4_VMS_L2D4PHI3Z1n2_wr_en;
wire [5:0] VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1_number;
wire [10:0] VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1;
VMStubs #("Tracklet") VMS_L2D4PHI3Z1n2(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z1n2),
.enable(VMR_L2D4_VMS_L2D4PHI3Z1n2_wr_en),
.number_out(VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1_number),
.read_add(VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1_read_add),
.data_out(VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z1n6;
wire VMR_L1D3_VMS_L1D3PHI3Z1n6_wr_en;
wire [5:0] VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1_number;
wire [10:0] VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1_read_add;
wire [17:0] VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1;
VMStubs #("Tracklet") VMS_L1D3PHI3Z1n6(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z1n6),
.enable(VMR_L1D3_VMS_L1D3PHI3Z1n6_wr_en),
.number_out(VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1_number),
.read_add(VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1_read_add),
.data_out(VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI4Z1n1;
wire VMR_L2D4_VMS_L2D4PHI4Z1n1_wr_en;
wire [5:0] VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1_number;
wire [10:0] VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1_read_add;
wire [17:0] VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1;
VMStubs #("Tracklet") VMS_L2D4PHI4Z1n1(
.data_in(VMR_L2D4_VMS_L2D4PHI4Z1n1),
.enable(VMR_L2D4_VMS_L2D4PHI4Z1n1_wr_en),
.number_out(VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1_number),
.read_add(VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1_read_add),
.data_out(VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z2n3;
wire VMR_L1D3_VMS_L1D3PHI1Z2n3_wr_en;
wire [5:0] VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1_number;
wire [10:0] VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1_read_add;
wire [17:0] VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1;
VMStubs #("Tracklet") VMS_L1D3PHI1Z2n3(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z2n3),
.enable(VMR_L1D3_VMS_L1D3PHI1Z2n3_wr_en),
.number_out(VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1_number),
.read_add(VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1_read_add),
.data_out(VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI1Z1n2;
wire VMR_L2D4_VMS_L2D4PHI1Z1n2_wr_en;
wire [5:0] VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1_number;
wire [10:0] VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1_read_add;
wire [17:0] VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1;
VMStubs #("Tracklet") VMS_L2D4PHI1Z1n2(
.data_in(VMR_L2D4_VMS_L2D4PHI1Z1n2),
.enable(VMR_L2D4_VMS_L2D4PHI1Z1n2_wr_en),
.number_out(VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1_number),
.read_add(VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1_read_add),
.data_out(VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z2n4;
wire VMR_L1D3_VMS_L1D3PHI1Z2n4_wr_en;
wire [5:0] VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1_number;
wire [10:0] VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1;
VMStubs #("Tracklet") VMS_L1D3PHI1Z2n4(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z2n4),
.enable(VMR_L1D3_VMS_L1D3PHI1Z2n4_wr_en),
.number_out(VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1_number),
.read_add(VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1_read_add),
.data_out(VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z1n3;
wire VMR_L2D4_VMS_L2D4PHI2Z1n3_wr_en;
wire [5:0] VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1_number;
wire [10:0] VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1;
VMStubs #("Tracklet") VMS_L2D4PHI2Z1n3(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z1n3),
.enable(VMR_L2D4_VMS_L2D4PHI2Z1n3_wr_en),
.number_out(VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1_number),
.read_add(VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1_read_add),
.data_out(VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z2n3;
wire VMR_L1D3_VMS_L1D3PHI2Z2n3_wr_en;
wire [5:0] VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1_number;
wire [10:0] VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1;
VMStubs #("Tracklet") VMS_L1D3PHI2Z2n3(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z2n3),
.enable(VMR_L1D3_VMS_L1D3PHI2Z2n3_wr_en),
.number_out(VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1_number),
.read_add(VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1_read_add),
.data_out(VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z1n4;
wire VMR_L2D4_VMS_L2D4PHI2Z1n4_wr_en;
wire [5:0] VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1_number;
wire [10:0] VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1;
VMStubs #("Tracklet") VMS_L2D4PHI2Z1n4(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z1n4),
.enable(VMR_L2D4_VMS_L2D4PHI2Z1n4_wr_en),
.number_out(VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1_number),
.read_add(VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1_read_add),
.data_out(VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z2n4;
wire VMR_L1D3_VMS_L1D3PHI2Z2n4_wr_en;
wire [5:0] VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1_number;
wire [10:0] VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1;
VMStubs #("Tracklet") VMS_L1D3PHI2Z2n4(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z2n4),
.enable(VMR_L1D3_VMS_L1D3PHI2Z2n4_wr_en),
.number_out(VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1_number),
.read_add(VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1_read_add),
.data_out(VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z1n3;
wire VMR_L2D4_VMS_L2D4PHI3Z1n3_wr_en;
wire [5:0] VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1_number;
wire [10:0] VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1;
VMStubs #("Tracklet") VMS_L2D4PHI3Z1n3(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z1n3),
.enable(VMR_L2D4_VMS_L2D4PHI3Z1n3_wr_en),
.number_out(VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1_number),
.read_add(VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1_read_add),
.data_out(VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z2n3;
wire VMR_L1D3_VMS_L1D3PHI3Z2n3_wr_en;
wire [5:0] VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1_number;
wire [10:0] VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1;
VMStubs #("Tracklet") VMS_L1D3PHI3Z2n3(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z2n3),
.enable(VMR_L1D3_VMS_L1D3PHI3Z2n3_wr_en),
.number_out(VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1_number),
.read_add(VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1_read_add),
.data_out(VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z1n4;
wire VMR_L2D4_VMS_L2D4PHI3Z1n4_wr_en;
wire [5:0] VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1_number;
wire [10:0] VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1;
VMStubs #("Tracklet") VMS_L2D4PHI3Z1n4(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z1n4),
.enable(VMR_L2D4_VMS_L2D4PHI3Z1n4_wr_en),
.number_out(VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1_number),
.read_add(VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1_read_add),
.data_out(VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z2n4;
wire VMR_L1D3_VMS_L1D3PHI3Z2n4_wr_en;
wire [5:0] VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1_number;
wire [10:0] VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1_read_add;
wire [17:0] VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1;
VMStubs #("Tracklet") VMS_L1D3PHI3Z2n4(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z2n4),
.enable(VMR_L1D3_VMS_L1D3PHI3Z2n4_wr_en),
.number_out(VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1_number),
.read_add(VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1_read_add),
.data_out(VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI4Z1n2;
wire VMR_L2D4_VMS_L2D4PHI4Z1n2_wr_en;
wire [5:0] VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1_number;
wire [10:0] VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1_read_add;
wire [17:0] VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1;
VMStubs #("Tracklet") VMS_L2D4PHI4Z1n2(
.data_in(VMR_L2D4_VMS_L2D4PHI4Z1n2),
.enable(VMR_L2D4_VMS_L2D4PHI4Z1n2_wr_en),
.number_out(VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1_number),
.read_add(VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1_read_add),
.data_out(VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z2n5;
wire VMR_L1D3_VMS_L1D3PHI1Z2n5_wr_en;
wire [5:0] VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2_number;
wire [10:0] VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2_read_add;
wire [17:0] VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2;
VMStubs #("Tracklet") VMS_L1D3PHI1Z2n5(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z2n5),
.enable(VMR_L1D3_VMS_L1D3PHI1Z2n5_wr_en),
.number_out(VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2_number),
.read_add(VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2_read_add),
.data_out(VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI1Z2n1;
wire VMR_L2D4_VMS_L2D4PHI1Z2n1_wr_en;
wire [5:0] VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2_number;
wire [10:0] VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2_read_add;
wire [17:0] VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2;
VMStubs #("Tracklet") VMS_L2D4PHI1Z2n1(
.data_in(VMR_L2D4_VMS_L2D4PHI1Z2n1),
.enable(VMR_L2D4_VMS_L2D4PHI1Z2n1_wr_en),
.number_out(VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2_number),
.read_add(VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2_read_add),
.data_out(VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z2n6;
wire VMR_L1D3_VMS_L1D3PHI1Z2n6_wr_en;
wire [5:0] VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2_number;
wire [10:0] VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2;
VMStubs #("Tracklet") VMS_L1D3PHI1Z2n6(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z2n6),
.enable(VMR_L1D3_VMS_L1D3PHI1Z2n6_wr_en),
.number_out(VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2_number),
.read_add(VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2_read_add),
.data_out(VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z2n1;
wire VMR_L2D4_VMS_L2D4PHI2Z2n1_wr_en;
wire [5:0] VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2_number;
wire [10:0] VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2;
VMStubs #("Tracklet") VMS_L2D4PHI2Z2n1(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z2n1),
.enable(VMR_L2D4_VMS_L2D4PHI2Z2n1_wr_en),
.number_out(VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2_number),
.read_add(VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2_read_add),
.data_out(VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z2n5;
wire VMR_L1D3_VMS_L1D3PHI2Z2n5_wr_en;
wire [5:0] VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2_number;
wire [10:0] VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2;
VMStubs #("Tracklet") VMS_L1D3PHI2Z2n5(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z2n5),
.enable(VMR_L1D3_VMS_L1D3PHI2Z2n5_wr_en),
.number_out(VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2_number),
.read_add(VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2_read_add),
.data_out(VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z2n2;
wire VMR_L2D4_VMS_L2D4PHI2Z2n2_wr_en;
wire [5:0] VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2_number;
wire [10:0] VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2;
VMStubs #("Tracklet") VMS_L2D4PHI2Z2n2(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z2n2),
.enable(VMR_L2D4_VMS_L2D4PHI2Z2n2_wr_en),
.number_out(VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2_number),
.read_add(VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2_read_add),
.data_out(VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z2n6;
wire VMR_L1D3_VMS_L1D3PHI2Z2n6_wr_en;
wire [5:0] VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2_number;
wire [10:0] VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2;
VMStubs #("Tracklet") VMS_L1D3PHI2Z2n6(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z2n6),
.enable(VMR_L1D3_VMS_L1D3PHI2Z2n6_wr_en),
.number_out(VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2_number),
.read_add(VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2_read_add),
.data_out(VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z2n1;
wire VMR_L2D4_VMS_L2D4PHI3Z2n1_wr_en;
wire [5:0] VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2_number;
wire [10:0] VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2;
VMStubs #("Tracklet") VMS_L2D4PHI3Z2n1(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z2n1),
.enable(VMR_L2D4_VMS_L2D4PHI3Z2n1_wr_en),
.number_out(VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2_number),
.read_add(VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2_read_add),
.data_out(VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z2n5;
wire VMR_L1D3_VMS_L1D3PHI3Z2n5_wr_en;
wire [5:0] VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2_number;
wire [10:0] VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2;
VMStubs #("Tracklet") VMS_L1D3PHI3Z2n5(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z2n5),
.enable(VMR_L1D3_VMS_L1D3PHI3Z2n5_wr_en),
.number_out(VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2_number),
.read_add(VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2_read_add),
.data_out(VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z2n2;
wire VMR_L2D4_VMS_L2D4PHI3Z2n2_wr_en;
wire [5:0] VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2_number;
wire [10:0] VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2;
VMStubs #("Tracklet") VMS_L2D4PHI3Z2n2(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z2n2),
.enable(VMR_L2D4_VMS_L2D4PHI3Z2n2_wr_en),
.number_out(VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2_number),
.read_add(VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2_read_add),
.data_out(VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z2n6;
wire VMR_L1D3_VMS_L1D3PHI3Z2n6_wr_en;
wire [5:0] VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2_number;
wire [10:0] VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2_read_add;
wire [17:0] VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2;
VMStubs #("Tracklet") VMS_L1D3PHI3Z2n6(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z2n6),
.enable(VMR_L1D3_VMS_L1D3PHI3Z2n6_wr_en),
.number_out(VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2_number),
.read_add(VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2_read_add),
.data_out(VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI4Z2n1;
wire VMR_L2D4_VMS_L2D4PHI4Z2n1_wr_en;
wire [5:0] VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2_number;
wire [10:0] VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2_read_add;
wire [17:0] VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2;
VMStubs #("Tracklet") VMS_L2D4PHI4Z2n1(
.data_in(VMR_L2D4_VMS_L2D4PHI4Z2n1),
.enable(VMR_L2D4_VMS_L2D4PHI4Z2n1_wr_en),
.number_out(VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2_number),
.read_add(VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2_read_add),
.data_out(VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI1Z1n1;
wire VMR_L1D4_VMS_L1D4PHI1Z1n1_wr_en;
wire [5:0] VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2_number;
wire [10:0] VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2_read_add;
wire [17:0] VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2;
VMStubs #("Tracklet") VMS_L1D4PHI1Z1n1(
.data_in(VMR_L1D4_VMS_L1D4PHI1Z1n1),
.enable(VMR_L1D4_VMS_L1D4PHI1Z1n1_wr_en),
.number_out(VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2_number),
.read_add(VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2_read_add),
.data_out(VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI1Z2n2;
wire VMR_L2D4_VMS_L2D4PHI1Z2n2_wr_en;
wire [5:0] VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2_number;
wire [10:0] VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2_read_add;
wire [17:0] VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2;
VMStubs #("Tracklet") VMS_L2D4PHI1Z2n2(
.data_in(VMR_L2D4_VMS_L2D4PHI1Z2n2),
.enable(VMR_L2D4_VMS_L2D4PHI1Z2n2_wr_en),
.number_out(VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2_number),
.read_add(VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2_read_add),
.data_out(VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI1Z1n2;
wire VMR_L1D4_VMS_L1D4PHI1Z1n2_wr_en;
wire [5:0] VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2_number;
wire [10:0] VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2;
VMStubs #("Tracklet") VMS_L1D4PHI1Z1n2(
.data_in(VMR_L1D4_VMS_L1D4PHI1Z1n2),
.enable(VMR_L1D4_VMS_L1D4PHI1Z1n2_wr_en),
.number_out(VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2_number),
.read_add(VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2_read_add),
.data_out(VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z2n3;
wire VMR_L2D4_VMS_L2D4PHI2Z2n3_wr_en;
wire [5:0] VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2_number;
wire [10:0] VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2;
VMStubs #("Tracklet") VMS_L2D4PHI2Z2n3(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z2n3),
.enable(VMR_L2D4_VMS_L2D4PHI2Z2n3_wr_en),
.number_out(VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2_number),
.read_add(VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2_read_add),
.data_out(VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI2Z1n1;
wire VMR_L1D4_VMS_L1D4PHI2Z1n1_wr_en;
wire [5:0] VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2_number;
wire [10:0] VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2;
VMStubs #("Tracklet") VMS_L1D4PHI2Z1n1(
.data_in(VMR_L1D4_VMS_L1D4PHI2Z1n1),
.enable(VMR_L1D4_VMS_L1D4PHI2Z1n1_wr_en),
.number_out(VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2_number),
.read_add(VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2_read_add),
.data_out(VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z2n4;
wire VMR_L2D4_VMS_L2D4PHI2Z2n4_wr_en;
wire [5:0] VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2_number;
wire [10:0] VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2;
VMStubs #("Tracklet") VMS_L2D4PHI2Z2n4(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z2n4),
.enable(VMR_L2D4_VMS_L2D4PHI2Z2n4_wr_en),
.number_out(VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2_number),
.read_add(VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2_read_add),
.data_out(VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI2Z1n2;
wire VMR_L1D4_VMS_L1D4PHI2Z1n2_wr_en;
wire [5:0] VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2_number;
wire [10:0] VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2;
VMStubs #("Tracklet") VMS_L1D4PHI2Z1n2(
.data_in(VMR_L1D4_VMS_L1D4PHI2Z1n2),
.enable(VMR_L1D4_VMS_L1D4PHI2Z1n2_wr_en),
.number_out(VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2_number),
.read_add(VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2_read_add),
.data_out(VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z2n3;
wire VMR_L2D4_VMS_L2D4PHI3Z2n3_wr_en;
wire [5:0] VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2_number;
wire [10:0] VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2;
VMStubs #("Tracklet") VMS_L2D4PHI3Z2n3(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z2n3),
.enable(VMR_L2D4_VMS_L2D4PHI3Z2n3_wr_en),
.number_out(VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2_number),
.read_add(VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2_read_add),
.data_out(VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI3Z1n1;
wire VMR_L1D4_VMS_L1D4PHI3Z1n1_wr_en;
wire [5:0] VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2_number;
wire [10:0] VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2;
VMStubs #("Tracklet") VMS_L1D4PHI3Z1n1(
.data_in(VMR_L1D4_VMS_L1D4PHI3Z1n1),
.enable(VMR_L1D4_VMS_L1D4PHI3Z1n1_wr_en),
.number_out(VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2_number),
.read_add(VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2_read_add),
.data_out(VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z2n4;
wire VMR_L2D4_VMS_L2D4PHI3Z2n4_wr_en;
wire [5:0] VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2_number;
wire [10:0] VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2;
VMStubs #("Tracklet") VMS_L2D4PHI3Z2n4(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z2n4),
.enable(VMR_L2D4_VMS_L2D4PHI3Z2n4_wr_en),
.number_out(VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2_number),
.read_add(VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2_read_add),
.data_out(VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI3Z1n2;
wire VMR_L1D4_VMS_L1D4PHI3Z1n2_wr_en;
wire [5:0] VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_number;
wire [10:0] VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_read_add;
wire [17:0] VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2;
VMStubs #("Tracklet") VMS_L1D4PHI3Z1n2(
.data_in(VMR_L1D4_VMS_L1D4PHI3Z1n2),
.enable(VMR_L1D4_VMS_L1D4PHI3Z1n2_wr_en),
.number_out(VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_number),
.read_add(VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_read_add),
.data_out(VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI4Z2n2;
wire VMR_L2D4_VMS_L2D4PHI4Z2n2_wr_en;
wire [5:0] VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_number;
wire [10:0] VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_read_add;
wire [17:0] VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2;
VMStubs #("Tracklet") VMS_L2D4PHI4Z2n2(
.data_in(VMR_L2D4_VMS_L2D4PHI4Z2n2),
.enable(VMR_L2D4_VMS_L2D4PHI4Z2n2_wr_en),
.number_out(VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_number),
.read_add(VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_read_add),
.data_out(VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z1n1;
wire VMR_L3D3_VMS_L3D3PHI1Z1n1_wr_en;
wire [5:0] VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_number;
wire [10:0] VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_read_add;
wire [17:0] VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1;
VMStubs #("Tracklet") VMS_L3D3PHI1Z1n1(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z1n1),
.enable(VMR_L3D3_VMS_L3D3PHI1Z1n1_wr_en),
.number_out(VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_number),
.read_add(VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_read_add),
.data_out(VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI1Z1n1;
wire VMR_L4D3_VMS_L4D3PHI1Z1n1_wr_en;
wire [5:0] VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_number;
wire [10:0] VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_read_add;
wire [17:0] VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1;
VMStubs #("Tracklet") VMS_L4D3PHI1Z1n1(
.data_in(VMR_L4D3_VMS_L4D3PHI1Z1n1),
.enable(VMR_L4D3_VMS_L4D3PHI1Z1n1_wr_en),
.number_out(VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_number),
.read_add(VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_read_add),
.data_out(VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z1n2;
wire VMR_L3D3_VMS_L3D3PHI1Z1n2_wr_en;
wire [5:0] VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1_number;
wire [10:0] VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1_read_add;
wire [17:0] VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1;
VMStubs #("Tracklet") VMS_L3D3PHI1Z1n2(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z1n2),
.enable(VMR_L3D3_VMS_L3D3PHI1Z1n2_wr_en),
.number_out(VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1_number),
.read_add(VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1_read_add),
.data_out(VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z1n1;
wire VMR_L4D3_VMS_L4D3PHI2Z1n1_wr_en;
wire [5:0] VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1_number;
wire [10:0] VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1_read_add;
wire [17:0] VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1;
VMStubs #("Tracklet") VMS_L4D3PHI2Z1n1(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z1n1),
.enable(VMR_L4D3_VMS_L4D3PHI2Z1n1_wr_en),
.number_out(VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1_number),
.read_add(VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1_read_add),
.data_out(VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z1n1;
wire VMR_L3D3_VMS_L3D3PHI2Z1n1_wr_en;
wire [5:0] VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1_number;
wire [10:0] VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1_read_add;
wire [17:0] VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1;
VMStubs #("Tracklet") VMS_L3D3PHI2Z1n1(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z1n1),
.enable(VMR_L3D3_VMS_L3D3PHI2Z1n1_wr_en),
.number_out(VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1_number),
.read_add(VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1_read_add),
.data_out(VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z1n2;
wire VMR_L4D3_VMS_L4D3PHI2Z1n2_wr_en;
wire [5:0] VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1_number;
wire [10:0] VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1_read_add;
wire [17:0] VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1;
VMStubs #("Tracklet") VMS_L4D3PHI2Z1n2(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z1n2),
.enable(VMR_L4D3_VMS_L4D3PHI2Z1n2_wr_en),
.number_out(VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1_number),
.read_add(VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1_read_add),
.data_out(VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z1n2;
wire VMR_L3D3_VMS_L3D3PHI2Z1n2_wr_en;
wire [5:0] VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1_number;
wire [10:0] VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1_read_add;
wire [17:0] VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1;
VMStubs #("Tracklet") VMS_L3D3PHI2Z1n2(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z1n2),
.enable(VMR_L3D3_VMS_L3D3PHI2Z1n2_wr_en),
.number_out(VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1_number),
.read_add(VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1_read_add),
.data_out(VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z1n1;
wire VMR_L4D3_VMS_L4D3PHI3Z1n1_wr_en;
wire [5:0] VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1_number;
wire [10:0] VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1_read_add;
wire [17:0] VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1;
VMStubs #("Tracklet") VMS_L4D3PHI3Z1n1(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z1n1),
.enable(VMR_L4D3_VMS_L4D3PHI3Z1n1_wr_en),
.number_out(VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1_number),
.read_add(VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1_read_add),
.data_out(VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z1n1;
wire VMR_L3D3_VMS_L3D3PHI3Z1n1_wr_en;
wire [5:0] VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1_number;
wire [10:0] VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1_read_add;
wire [17:0] VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1;
VMStubs #("Tracklet") VMS_L3D3PHI3Z1n1(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z1n1),
.enable(VMR_L3D3_VMS_L3D3PHI3Z1n1_wr_en),
.number_out(VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1_number),
.read_add(VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1_read_add),
.data_out(VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z1n2;
wire VMR_L4D3_VMS_L4D3PHI3Z1n2_wr_en;
wire [5:0] VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1_number;
wire [10:0] VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1_read_add;
wire [17:0] VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1;
VMStubs #("Tracklet") VMS_L4D3PHI3Z1n2(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z1n2),
.enable(VMR_L4D3_VMS_L4D3PHI3Z1n2_wr_en),
.number_out(VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1_number),
.read_add(VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1_read_add),
.data_out(VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z1n2;
wire VMR_L3D3_VMS_L3D3PHI3Z1n2_wr_en;
wire [5:0] VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1_number;
wire [10:0] VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1_read_add;
wire [17:0] VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1;
VMStubs #("Tracklet") VMS_L3D3PHI3Z1n2(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z1n2),
.enable(VMR_L3D3_VMS_L3D3PHI3Z1n2_wr_en),
.number_out(VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1_number),
.read_add(VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1_read_add),
.data_out(VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI4Z1n1;
wire VMR_L4D3_VMS_L4D3PHI4Z1n1_wr_en;
wire [5:0] VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1_number;
wire [10:0] VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1_read_add;
wire [17:0] VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1;
VMStubs #("Tracklet") VMS_L4D3PHI4Z1n1(
.data_in(VMR_L4D3_VMS_L4D3PHI4Z1n1),
.enable(VMR_L4D3_VMS_L4D3PHI4Z1n1_wr_en),
.number_out(VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1_number),
.read_add(VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1_read_add),
.data_out(VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z2n1;
wire VMR_L3D3_VMS_L3D3PHI1Z2n1_wr_en;
wire [5:0] VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_number;
wire [10:0] VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_read_add;
wire [17:0] VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2;
VMStubs #("Tracklet") VMS_L3D3PHI1Z2n1(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z2n1),
.enable(VMR_L3D3_VMS_L3D3PHI1Z2n1_wr_en),
.number_out(VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_number),
.read_add(VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_read_add),
.data_out(VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI1Z2n1;
wire VMR_L4D3_VMS_L4D3PHI1Z2n1_wr_en;
wire [5:0] VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_number;
wire [10:0] VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_read_add;
wire [17:0] VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2;
VMStubs #("Tracklet") VMS_L4D3PHI1Z2n1(
.data_in(VMR_L4D3_VMS_L4D3PHI1Z2n1),
.enable(VMR_L4D3_VMS_L4D3PHI1Z2n1_wr_en),
.number_out(VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_number),
.read_add(VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_read_add),
.data_out(VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z2n2;
wire VMR_L3D3_VMS_L3D3PHI1Z2n2_wr_en;
wire [5:0] VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2_number;
wire [10:0] VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2;
VMStubs #("Tracklet") VMS_L3D3PHI1Z2n2(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z2n2),
.enable(VMR_L3D3_VMS_L3D3PHI1Z2n2_wr_en),
.number_out(VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2_number),
.read_add(VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2_read_add),
.data_out(VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z2n1;
wire VMR_L4D3_VMS_L4D3PHI2Z2n1_wr_en;
wire [5:0] VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2_number;
wire [10:0] VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2;
VMStubs #("Tracklet") VMS_L4D3PHI2Z2n1(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z2n1),
.enable(VMR_L4D3_VMS_L4D3PHI2Z2n1_wr_en),
.number_out(VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2_number),
.read_add(VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2_read_add),
.data_out(VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z2n1;
wire VMR_L3D3_VMS_L3D3PHI2Z2n1_wr_en;
wire [5:0] VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2_number;
wire [10:0] VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2;
VMStubs #("Tracklet") VMS_L3D3PHI2Z2n1(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z2n1),
.enable(VMR_L3D3_VMS_L3D3PHI2Z2n1_wr_en),
.number_out(VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2_number),
.read_add(VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2_read_add),
.data_out(VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z2n2;
wire VMR_L4D3_VMS_L4D3PHI2Z2n2_wr_en;
wire [5:0] VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2_number;
wire [10:0] VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2;
VMStubs #("Tracklet") VMS_L4D3PHI2Z2n2(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z2n2),
.enable(VMR_L4D3_VMS_L4D3PHI2Z2n2_wr_en),
.number_out(VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2_number),
.read_add(VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2_read_add),
.data_out(VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z2n2;
wire VMR_L3D3_VMS_L3D3PHI2Z2n2_wr_en;
wire [5:0] VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2_number;
wire [10:0] VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2;
VMStubs #("Tracklet") VMS_L3D3PHI2Z2n2(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z2n2),
.enable(VMR_L3D3_VMS_L3D3PHI2Z2n2_wr_en),
.number_out(VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2_number),
.read_add(VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2_read_add),
.data_out(VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z2n1;
wire VMR_L4D3_VMS_L4D3PHI3Z2n1_wr_en;
wire [5:0] VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2_number;
wire [10:0] VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2;
VMStubs #("Tracklet") VMS_L4D3PHI3Z2n1(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z2n1),
.enable(VMR_L4D3_VMS_L4D3PHI3Z2n1_wr_en),
.number_out(VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2_number),
.read_add(VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2_read_add),
.data_out(VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z2n1;
wire VMR_L3D3_VMS_L3D3PHI3Z2n1_wr_en;
wire [5:0] VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2_number;
wire [10:0] VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2;
VMStubs #("Tracklet") VMS_L3D3PHI3Z2n1(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z2n1),
.enable(VMR_L3D3_VMS_L3D3PHI3Z2n1_wr_en),
.number_out(VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2_number),
.read_add(VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2_read_add),
.data_out(VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z2n2;
wire VMR_L4D3_VMS_L4D3PHI3Z2n2_wr_en;
wire [5:0] VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2_number;
wire [10:0] VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2;
VMStubs #("Tracklet") VMS_L4D3PHI3Z2n2(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z2n2),
.enable(VMR_L4D3_VMS_L4D3PHI3Z2n2_wr_en),
.number_out(VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2_number),
.read_add(VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2_read_add),
.data_out(VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z2n2;
wire VMR_L3D3_VMS_L3D3PHI3Z2n2_wr_en;
wire [5:0] VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2_number;
wire [10:0] VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2_read_add;
wire [17:0] VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2;
VMStubs #("Tracklet") VMS_L3D3PHI3Z2n2(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z2n2),
.enable(VMR_L3D3_VMS_L3D3PHI3Z2n2_wr_en),
.number_out(VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2_number),
.read_add(VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2_read_add),
.data_out(VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI4Z2n1;
wire VMR_L4D3_VMS_L4D3PHI4Z2n1_wr_en;
wire [5:0] VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2_number;
wire [10:0] VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2_read_add;
wire [17:0] VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2;
VMStubs #("Tracklet") VMS_L4D3PHI4Z2n1(
.data_in(VMR_L4D3_VMS_L4D3PHI4Z2n1),
.enable(VMR_L4D3_VMS_L4D3PHI4Z2n1_wr_en),
.number_out(VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2_number),
.read_add(VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2_read_add),
.data_out(VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z1n3;
wire VMR_L3D3_VMS_L3D3PHI1Z1n3_wr_en;
wire [5:0] VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2_number;
wire [10:0] VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2_read_add;
wire [17:0] VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2;
VMStubs #("Tracklet") VMS_L3D3PHI1Z1n3(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z1n3),
.enable(VMR_L3D3_VMS_L3D3PHI1Z1n3_wr_en),
.number_out(VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2_number),
.read_add(VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2_read_add),
.data_out(VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI1Z2n2;
wire VMR_L4D3_VMS_L4D3PHI1Z2n2_wr_en;
wire [5:0] VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2_number;
wire [10:0] VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2_read_add;
wire [17:0] VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2;
VMStubs #("Tracklet") VMS_L4D3PHI1Z2n2(
.data_in(VMR_L4D3_VMS_L4D3PHI1Z2n2),
.enable(VMR_L4D3_VMS_L4D3PHI1Z2n2_wr_en),
.number_out(VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2_number),
.read_add(VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2_read_add),
.data_out(VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z1n4;
wire VMR_L3D3_VMS_L3D3PHI1Z1n4_wr_en;
wire [5:0] VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2_number;
wire [10:0] VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2;
VMStubs #("Tracklet") VMS_L3D3PHI1Z1n4(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z1n4),
.enable(VMR_L3D3_VMS_L3D3PHI1Z1n4_wr_en),
.number_out(VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2_number),
.read_add(VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2_read_add),
.data_out(VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z2n3;
wire VMR_L4D3_VMS_L4D3PHI2Z2n3_wr_en;
wire [5:0] VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2_number;
wire [10:0] VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2;
VMStubs #("Tracklet") VMS_L4D3PHI2Z2n3(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z2n3),
.enable(VMR_L4D3_VMS_L4D3PHI2Z2n3_wr_en),
.number_out(VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2_number),
.read_add(VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2_read_add),
.data_out(VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z1n3;
wire VMR_L3D3_VMS_L3D3PHI2Z1n3_wr_en;
wire [5:0] VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2_number;
wire [10:0] VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2;
VMStubs #("Tracklet") VMS_L3D3PHI2Z1n3(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z1n3),
.enable(VMR_L3D3_VMS_L3D3PHI2Z1n3_wr_en),
.number_out(VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2_number),
.read_add(VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2_read_add),
.data_out(VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z2n4;
wire VMR_L4D3_VMS_L4D3PHI2Z2n4_wr_en;
wire [5:0] VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2_number;
wire [10:0] VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2;
VMStubs #("Tracklet") VMS_L4D3PHI2Z2n4(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z2n4),
.enable(VMR_L4D3_VMS_L4D3PHI2Z2n4_wr_en),
.number_out(VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2_number),
.read_add(VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2_read_add),
.data_out(VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z1n4;
wire VMR_L3D3_VMS_L3D3PHI2Z1n4_wr_en;
wire [5:0] VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2_number;
wire [10:0] VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2;
VMStubs #("Tracklet") VMS_L3D3PHI2Z1n4(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z1n4),
.enable(VMR_L3D3_VMS_L3D3PHI2Z1n4_wr_en),
.number_out(VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2_number),
.read_add(VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2_read_add),
.data_out(VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z2n3;
wire VMR_L4D3_VMS_L4D3PHI3Z2n3_wr_en;
wire [5:0] VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2_number;
wire [10:0] VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2;
VMStubs #("Tracklet") VMS_L4D3PHI3Z2n3(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z2n3),
.enable(VMR_L4D3_VMS_L4D3PHI3Z2n3_wr_en),
.number_out(VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2_number),
.read_add(VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2_read_add),
.data_out(VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z1n3;
wire VMR_L3D3_VMS_L3D3PHI3Z1n3_wr_en;
wire [5:0] VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2_number;
wire [10:0] VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2;
VMStubs #("Tracklet") VMS_L3D3PHI3Z1n3(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z1n3),
.enable(VMR_L3D3_VMS_L3D3PHI3Z1n3_wr_en),
.number_out(VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2_number),
.read_add(VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2_read_add),
.data_out(VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z2n4;
wire VMR_L4D3_VMS_L4D3PHI3Z2n4_wr_en;
wire [5:0] VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2_number;
wire [10:0] VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2;
VMStubs #("Tracklet") VMS_L4D3PHI3Z2n4(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z2n4),
.enable(VMR_L4D3_VMS_L4D3PHI3Z2n4_wr_en),
.number_out(VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2_number),
.read_add(VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2_read_add),
.data_out(VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z1n4;
wire VMR_L3D3_VMS_L3D3PHI3Z1n4_wr_en;
wire [5:0] VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2_number;
wire [10:0] VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2_read_add;
wire [17:0] VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2;
VMStubs #("Tracklet") VMS_L3D3PHI3Z1n4(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z1n4),
.enable(VMR_L3D3_VMS_L3D3PHI3Z1n4_wr_en),
.number_out(VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2_number),
.read_add(VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2_read_add),
.data_out(VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI4Z2n2;
wire VMR_L4D3_VMS_L4D3PHI4Z2n2_wr_en;
wire [5:0] VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2_number;
wire [10:0] VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2_read_add;
wire [17:0] VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2;
VMStubs #("Tracklet") VMS_L4D3PHI4Z2n2(
.data_in(VMR_L4D3_VMS_L4D3PHI4Z2n2),
.enable(VMR_L4D3_VMS_L4D3PHI4Z2n2_wr_en),
.number_out(VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2_number),
.read_add(VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2_read_add),
.data_out(VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z2n3;
wire VMR_L3D3_VMS_L3D3PHI1Z2n3_wr_en;
wire [5:0] VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1_number;
wire [10:0] VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1_read_add;
wire [17:0] VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1;
VMStubs #("Tracklet") VMS_L3D3PHI1Z2n3(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z2n3),
.enable(VMR_L3D3_VMS_L3D3PHI1Z2n3_wr_en),
.number_out(VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1_number),
.read_add(VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1_read_add),
.data_out(VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI1Z1n1;
wire VMR_L4D4_VMS_L4D4PHI1Z1n1_wr_en;
wire [5:0] VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1_number;
wire [10:0] VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1_read_add;
wire [17:0] VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1;
VMStubs #("Tracklet") VMS_L4D4PHI1Z1n1(
.data_in(VMR_L4D4_VMS_L4D4PHI1Z1n1),
.enable(VMR_L4D4_VMS_L4D4PHI1Z1n1_wr_en),
.number_out(VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1_number),
.read_add(VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1_read_add),
.data_out(VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z2n4;
wire VMR_L3D3_VMS_L3D3PHI1Z2n4_wr_en;
wire [5:0] VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1_number;
wire [10:0] VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1;
VMStubs #("Tracklet") VMS_L3D3PHI1Z2n4(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z2n4),
.enable(VMR_L3D3_VMS_L3D3PHI1Z2n4_wr_en),
.number_out(VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1_number),
.read_add(VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1_read_add),
.data_out(VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z1n1;
wire VMR_L4D4_VMS_L4D4PHI2Z1n1_wr_en;
wire [5:0] VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1_number;
wire [10:0] VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1;
VMStubs #("Tracklet") VMS_L4D4PHI2Z1n1(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z1n1),
.enable(VMR_L4D4_VMS_L4D4PHI2Z1n1_wr_en),
.number_out(VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1_number),
.read_add(VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1_read_add),
.data_out(VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z2n3;
wire VMR_L3D3_VMS_L3D3PHI2Z2n3_wr_en;
wire [5:0] VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1_number;
wire [10:0] VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1;
VMStubs #("Tracklet") VMS_L3D3PHI2Z2n3(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z2n3),
.enable(VMR_L3D3_VMS_L3D3PHI2Z2n3_wr_en),
.number_out(VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1_number),
.read_add(VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1_read_add),
.data_out(VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z1n2;
wire VMR_L4D4_VMS_L4D4PHI2Z1n2_wr_en;
wire [5:0] VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1_number;
wire [10:0] VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1;
VMStubs #("Tracklet") VMS_L4D4PHI2Z1n2(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z1n2),
.enable(VMR_L4D4_VMS_L4D4PHI2Z1n2_wr_en),
.number_out(VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1_number),
.read_add(VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1_read_add),
.data_out(VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z2n4;
wire VMR_L3D3_VMS_L3D3PHI2Z2n4_wr_en;
wire [5:0] VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1_number;
wire [10:0] VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1;
VMStubs #("Tracklet") VMS_L3D3PHI2Z2n4(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z2n4),
.enable(VMR_L3D3_VMS_L3D3PHI2Z2n4_wr_en),
.number_out(VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1_number),
.read_add(VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1_read_add),
.data_out(VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z1n1;
wire VMR_L4D4_VMS_L4D4PHI3Z1n1_wr_en;
wire [5:0] VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1_number;
wire [10:0] VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1;
VMStubs #("Tracklet") VMS_L4D4PHI3Z1n1(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z1n1),
.enable(VMR_L4D4_VMS_L4D4PHI3Z1n1_wr_en),
.number_out(VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1_number),
.read_add(VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1_read_add),
.data_out(VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z2n3;
wire VMR_L3D3_VMS_L3D3PHI3Z2n3_wr_en;
wire [5:0] VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1_number;
wire [10:0] VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1;
VMStubs #("Tracklet") VMS_L3D3PHI3Z2n3(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z2n3),
.enable(VMR_L3D3_VMS_L3D3PHI3Z2n3_wr_en),
.number_out(VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1_number),
.read_add(VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1_read_add),
.data_out(VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z1n2;
wire VMR_L4D4_VMS_L4D4PHI3Z1n2_wr_en;
wire [5:0] VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1_number;
wire [10:0] VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1;
VMStubs #("Tracklet") VMS_L4D4PHI3Z1n2(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z1n2),
.enable(VMR_L4D4_VMS_L4D4PHI3Z1n2_wr_en),
.number_out(VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1_number),
.read_add(VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1_read_add),
.data_out(VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z2n4;
wire VMR_L3D3_VMS_L3D3PHI3Z2n4_wr_en;
wire [5:0] VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1_number;
wire [10:0] VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1_read_add;
wire [17:0] VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1;
VMStubs #("Tracklet") VMS_L3D3PHI3Z2n4(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z2n4),
.enable(VMR_L3D3_VMS_L3D3PHI3Z2n4_wr_en),
.number_out(VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1_number),
.read_add(VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1_read_add),
.data_out(VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI4Z1n1;
wire VMR_L4D4_VMS_L4D4PHI4Z1n1_wr_en;
wire [5:0] VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1_number;
wire [10:0] VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1_read_add;
wire [17:0] VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1;
VMStubs #("Tracklet") VMS_L4D4PHI4Z1n1(
.data_in(VMR_L4D4_VMS_L4D4PHI4Z1n1),
.enable(VMR_L4D4_VMS_L4D4PHI4Z1n1_wr_en),
.number_out(VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1_number),
.read_add(VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1_read_add),
.data_out(VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z1n1;
wire VMR_L3D4_VMS_L3D4PHI1Z1n1_wr_en;
wire [5:0] VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1_number;
wire [10:0] VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1_read_add;
wire [17:0] VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1;
VMStubs #("Tracklet") VMS_L3D4PHI1Z1n1(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z1n1),
.enable(VMR_L3D4_VMS_L3D4PHI1Z1n1_wr_en),
.number_out(VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1_number),
.read_add(VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1_read_add),
.data_out(VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI1Z1n2;
wire VMR_L4D4_VMS_L4D4PHI1Z1n2_wr_en;
wire [5:0] VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1_number;
wire [10:0] VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1_read_add;
wire [17:0] VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1;
VMStubs #("Tracklet") VMS_L4D4PHI1Z1n2(
.data_in(VMR_L4D4_VMS_L4D4PHI1Z1n2),
.enable(VMR_L4D4_VMS_L4D4PHI1Z1n2_wr_en),
.number_out(VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1_number),
.read_add(VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1_read_add),
.data_out(VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z1n2;
wire VMR_L3D4_VMS_L3D4PHI1Z1n2_wr_en;
wire [5:0] VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1_number;
wire [10:0] VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1;
VMStubs #("Tracklet") VMS_L3D4PHI1Z1n2(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z1n2),
.enable(VMR_L3D4_VMS_L3D4PHI1Z1n2_wr_en),
.number_out(VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1_number),
.read_add(VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1_read_add),
.data_out(VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z1n3;
wire VMR_L4D4_VMS_L4D4PHI2Z1n3_wr_en;
wire [5:0] VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1_number;
wire [10:0] VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1;
VMStubs #("Tracklet") VMS_L4D4PHI2Z1n3(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z1n3),
.enable(VMR_L4D4_VMS_L4D4PHI2Z1n3_wr_en),
.number_out(VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1_number),
.read_add(VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1_read_add),
.data_out(VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z1n1;
wire VMR_L3D4_VMS_L3D4PHI2Z1n1_wr_en;
wire [5:0] VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1_number;
wire [10:0] VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1;
VMStubs #("Tracklet") VMS_L3D4PHI2Z1n1(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z1n1),
.enable(VMR_L3D4_VMS_L3D4PHI2Z1n1_wr_en),
.number_out(VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1_number),
.read_add(VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1_read_add),
.data_out(VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z1n4;
wire VMR_L4D4_VMS_L4D4PHI2Z1n4_wr_en;
wire [5:0] VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1_number;
wire [10:0] VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1;
VMStubs #("Tracklet") VMS_L4D4PHI2Z1n4(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z1n4),
.enable(VMR_L4D4_VMS_L4D4PHI2Z1n4_wr_en),
.number_out(VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1_number),
.read_add(VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1_read_add),
.data_out(VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z1n2;
wire VMR_L3D4_VMS_L3D4PHI2Z1n2_wr_en;
wire [5:0] VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1_number;
wire [10:0] VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1;
VMStubs #("Tracklet") VMS_L3D4PHI2Z1n2(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z1n2),
.enable(VMR_L3D4_VMS_L3D4PHI2Z1n2_wr_en),
.number_out(VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1_number),
.read_add(VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1_read_add),
.data_out(VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z1n3;
wire VMR_L4D4_VMS_L4D4PHI3Z1n3_wr_en;
wire [5:0] VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1_number;
wire [10:0] VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1;
VMStubs #("Tracklet") VMS_L4D4PHI3Z1n3(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z1n3),
.enable(VMR_L4D4_VMS_L4D4PHI3Z1n3_wr_en),
.number_out(VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1_number),
.read_add(VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1_read_add),
.data_out(VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z1n1;
wire VMR_L3D4_VMS_L3D4PHI3Z1n1_wr_en;
wire [5:0] VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1_number;
wire [10:0] VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1;
VMStubs #("Tracklet") VMS_L3D4PHI3Z1n1(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z1n1),
.enable(VMR_L3D4_VMS_L3D4PHI3Z1n1_wr_en),
.number_out(VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1_number),
.read_add(VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1_read_add),
.data_out(VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z1n4;
wire VMR_L4D4_VMS_L4D4PHI3Z1n4_wr_en;
wire [5:0] VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1_number;
wire [10:0] VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1;
VMStubs #("Tracklet") VMS_L4D4PHI3Z1n4(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z1n4),
.enable(VMR_L4D4_VMS_L4D4PHI3Z1n4_wr_en),
.number_out(VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1_number),
.read_add(VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1_read_add),
.data_out(VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z1n2;
wire VMR_L3D4_VMS_L3D4PHI3Z1n2_wr_en;
wire [5:0] VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_number;
wire [10:0] VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_read_add;
wire [17:0] VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1;
VMStubs #("Tracklet") VMS_L3D4PHI3Z1n2(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z1n2),
.enable(VMR_L3D4_VMS_L3D4PHI3Z1n2_wr_en),
.number_out(VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_number),
.read_add(VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_read_add),
.data_out(VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI4Z1n2;
wire VMR_L4D4_VMS_L4D4PHI4Z1n2_wr_en;
wire [5:0] VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_number;
wire [10:0] VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_read_add;
wire [17:0] VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1;
VMStubs #("Tracklet") VMS_L4D4PHI4Z1n2(
.data_in(VMR_L4D4_VMS_L4D4PHI4Z1n2),
.enable(VMR_L4D4_VMS_L4D4PHI4Z1n2_wr_en),
.number_out(VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_number),
.read_add(VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_read_add),
.data_out(VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z1n3;
wire VMR_L3D4_VMS_L3D4PHI1Z1n3_wr_en;
wire [5:0] VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2_number;
wire [10:0] VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2_read_add;
wire [17:0] VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2;
VMStubs #("Tracklet") VMS_L3D4PHI1Z1n3(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z1n3),
.enable(VMR_L3D4_VMS_L3D4PHI1Z1n3_wr_en),
.number_out(VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2_number),
.read_add(VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2_read_add),
.data_out(VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI1Z2n1;
wire VMR_L4D4_VMS_L4D4PHI1Z2n1_wr_en;
wire [5:0] VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2_number;
wire [10:0] VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2_read_add;
wire [17:0] VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2;
VMStubs #("Tracklet") VMS_L4D4PHI1Z2n1(
.data_in(VMR_L4D4_VMS_L4D4PHI1Z2n1),
.enable(VMR_L4D4_VMS_L4D4PHI1Z2n1_wr_en),
.number_out(VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2_number),
.read_add(VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2_read_add),
.data_out(VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z1n4;
wire VMR_L3D4_VMS_L3D4PHI1Z1n4_wr_en;
wire [5:0] VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2_number;
wire [10:0] VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2;
VMStubs #("Tracklet") VMS_L3D4PHI1Z1n4(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z1n4),
.enable(VMR_L3D4_VMS_L3D4PHI1Z1n4_wr_en),
.number_out(VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2_number),
.read_add(VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2_read_add),
.data_out(VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z2n1;
wire VMR_L4D4_VMS_L4D4PHI2Z2n1_wr_en;
wire [5:0] VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2_number;
wire [10:0] VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2;
VMStubs #("Tracklet") VMS_L4D4PHI2Z2n1(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z2n1),
.enable(VMR_L4D4_VMS_L4D4PHI2Z2n1_wr_en),
.number_out(VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2_number),
.read_add(VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2_read_add),
.data_out(VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z1n3;
wire VMR_L3D4_VMS_L3D4PHI2Z1n3_wr_en;
wire [5:0] VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2_number;
wire [10:0] VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2;
VMStubs #("Tracklet") VMS_L3D4PHI2Z1n3(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z1n3),
.enable(VMR_L3D4_VMS_L3D4PHI2Z1n3_wr_en),
.number_out(VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2_number),
.read_add(VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2_read_add),
.data_out(VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z2n2;
wire VMR_L4D4_VMS_L4D4PHI2Z2n2_wr_en;
wire [5:0] VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2_number;
wire [10:0] VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2;
VMStubs #("Tracklet") VMS_L4D4PHI2Z2n2(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z2n2),
.enable(VMR_L4D4_VMS_L4D4PHI2Z2n2_wr_en),
.number_out(VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2_number),
.read_add(VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2_read_add),
.data_out(VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z1n4;
wire VMR_L3D4_VMS_L3D4PHI2Z1n4_wr_en;
wire [5:0] VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2_number;
wire [10:0] VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2;
VMStubs #("Tracklet") VMS_L3D4PHI2Z1n4(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z1n4),
.enable(VMR_L3D4_VMS_L3D4PHI2Z1n4_wr_en),
.number_out(VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2_number),
.read_add(VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2_read_add),
.data_out(VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z2n1;
wire VMR_L4D4_VMS_L4D4PHI3Z2n1_wr_en;
wire [5:0] VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2_number;
wire [10:0] VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2;
VMStubs #("Tracklet") VMS_L4D4PHI3Z2n1(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z2n1),
.enable(VMR_L4D4_VMS_L4D4PHI3Z2n1_wr_en),
.number_out(VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2_number),
.read_add(VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2_read_add),
.data_out(VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z1n3;
wire VMR_L3D4_VMS_L3D4PHI3Z1n3_wr_en;
wire [5:0] VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2_number;
wire [10:0] VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2;
VMStubs #("Tracklet") VMS_L3D4PHI3Z1n3(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z1n3),
.enable(VMR_L3D4_VMS_L3D4PHI3Z1n3_wr_en),
.number_out(VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2_number),
.read_add(VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2_read_add),
.data_out(VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z2n2;
wire VMR_L4D4_VMS_L4D4PHI3Z2n2_wr_en;
wire [5:0] VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2_number;
wire [10:0] VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2;
VMStubs #("Tracklet") VMS_L4D4PHI3Z2n2(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z2n2),
.enable(VMR_L4D4_VMS_L4D4PHI3Z2n2_wr_en),
.number_out(VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2_number),
.read_add(VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2_read_add),
.data_out(VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z1n4;
wire VMR_L3D4_VMS_L3D4PHI3Z1n4_wr_en;
wire [5:0] VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2_number;
wire [10:0] VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2_read_add;
wire [17:0] VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2;
VMStubs #("Tracklet") VMS_L3D4PHI3Z1n4(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z1n4),
.enable(VMR_L3D4_VMS_L3D4PHI3Z1n4_wr_en),
.number_out(VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2_number),
.read_add(VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2_read_add),
.data_out(VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI4Z2n1;
wire VMR_L4D4_VMS_L4D4PHI4Z2n1_wr_en;
wire [5:0] VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2_number;
wire [10:0] VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2_read_add;
wire [17:0] VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2;
VMStubs #("Tracklet") VMS_L4D4PHI4Z2n1(
.data_in(VMR_L4D4_VMS_L4D4PHI4Z2n1),
.enable(VMR_L4D4_VMS_L4D4PHI4Z2n1_wr_en),
.number_out(VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2_number),
.read_add(VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2_read_add),
.data_out(VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z2n1;
wire VMR_L3D4_VMS_L3D4PHI1Z2n1_wr_en;
wire [5:0] VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2_number;
wire [10:0] VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2_read_add;
wire [17:0] VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2;
VMStubs #("Tracklet") VMS_L3D4PHI1Z2n1(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z2n1),
.enable(VMR_L3D4_VMS_L3D4PHI1Z2n1_wr_en),
.number_out(VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2_number),
.read_add(VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2_read_add),
.data_out(VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI1Z2n2;
wire VMR_L4D4_VMS_L4D4PHI1Z2n2_wr_en;
wire [5:0] VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2_number;
wire [10:0] VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2_read_add;
wire [17:0] VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2;
VMStubs #("Tracklet") VMS_L4D4PHI1Z2n2(
.data_in(VMR_L4D4_VMS_L4D4PHI1Z2n2),
.enable(VMR_L4D4_VMS_L4D4PHI1Z2n2_wr_en),
.number_out(VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2_number),
.read_add(VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2_read_add),
.data_out(VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z2n2;
wire VMR_L3D4_VMS_L3D4PHI1Z2n2_wr_en;
wire [5:0] VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2_number;
wire [10:0] VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2;
VMStubs #("Tracklet") VMS_L3D4PHI1Z2n2(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z2n2),
.enable(VMR_L3D4_VMS_L3D4PHI1Z2n2_wr_en),
.number_out(VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2_number),
.read_add(VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2_read_add),
.data_out(VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z2n3;
wire VMR_L4D4_VMS_L4D4PHI2Z2n3_wr_en;
wire [5:0] VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2_number;
wire [10:0] VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2;
VMStubs #("Tracklet") VMS_L4D4PHI2Z2n3(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z2n3),
.enable(VMR_L4D4_VMS_L4D4PHI2Z2n3_wr_en),
.number_out(VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2_number),
.read_add(VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2_read_add),
.data_out(VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z2n1;
wire VMR_L3D4_VMS_L3D4PHI2Z2n1_wr_en;
wire [5:0] VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2_number;
wire [10:0] VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2;
VMStubs #("Tracklet") VMS_L3D4PHI2Z2n1(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z2n1),
.enable(VMR_L3D4_VMS_L3D4PHI2Z2n1_wr_en),
.number_out(VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2_number),
.read_add(VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2_read_add),
.data_out(VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z2n4;
wire VMR_L4D4_VMS_L4D4PHI2Z2n4_wr_en;
wire [5:0] VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2_number;
wire [10:0] VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2;
VMStubs #("Tracklet") VMS_L4D4PHI2Z2n4(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z2n4),
.enable(VMR_L4D4_VMS_L4D4PHI2Z2n4_wr_en),
.number_out(VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2_number),
.read_add(VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2_read_add),
.data_out(VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z2n2;
wire VMR_L3D4_VMS_L3D4PHI2Z2n2_wr_en;
wire [5:0] VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2_number;
wire [10:0] VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2;
VMStubs #("Tracklet") VMS_L3D4PHI2Z2n2(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z2n2),
.enable(VMR_L3D4_VMS_L3D4PHI2Z2n2_wr_en),
.number_out(VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2_number),
.read_add(VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2_read_add),
.data_out(VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z2n3;
wire VMR_L4D4_VMS_L4D4PHI3Z2n3_wr_en;
wire [5:0] VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2_number;
wire [10:0] VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2;
VMStubs #("Tracklet") VMS_L4D4PHI3Z2n3(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z2n3),
.enable(VMR_L4D4_VMS_L4D4PHI3Z2n3_wr_en),
.number_out(VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2_number),
.read_add(VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2_read_add),
.data_out(VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z2n1;
wire VMR_L3D4_VMS_L3D4PHI3Z2n1_wr_en;
wire [5:0] VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2_number;
wire [10:0] VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2;
VMStubs #("Tracklet") VMS_L3D4PHI3Z2n1(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z2n1),
.enable(VMR_L3D4_VMS_L3D4PHI3Z2n1_wr_en),
.number_out(VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2_number),
.read_add(VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2_read_add),
.data_out(VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z2n4;
wire VMR_L4D4_VMS_L4D4PHI3Z2n4_wr_en;
wire [5:0] VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2_number;
wire [10:0] VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2;
VMStubs #("Tracklet") VMS_L4D4PHI3Z2n4(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z2n4),
.enable(VMR_L4D4_VMS_L4D4PHI3Z2n4_wr_en),
.number_out(VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2_number),
.read_add(VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2_read_add),
.data_out(VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z2n2;
wire VMR_L3D4_VMS_L3D4PHI3Z2n2_wr_en;
wire [5:0] VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_number;
wire [10:0] VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_read_add;
wire [17:0] VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2;
VMStubs #("Tracklet") VMS_L3D4PHI3Z2n2(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z2n2),
.enable(VMR_L3D4_VMS_L3D4PHI3Z2n2_wr_en),
.number_out(VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_number),
.read_add(VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_read_add),
.data_out(VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI4Z2n2;
wire VMR_L4D4_VMS_L4D4PHI4Z2n2_wr_en;
wire [5:0] VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_number;
wire [10:0] VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_read_add;
wire [17:0] VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2;
VMStubs #("Tracklet") VMS_L4D4PHI4Z2n2(
.data_in(VMR_L4D4_VMS_L4D4PHI4Z2n2),
.enable(VMR_L4D4_VMS_L4D4PHI4Z2n2_wr_en),
.number_out(VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_number),
.read_add(VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_read_add),
.data_out(VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z1n1;
wire VMR_L5D3_VMS_L5D3PHI1Z1n1_wr_en;
wire [5:0] VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_number;
wire [10:0] VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_read_add;
wire [17:0] VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1;
VMStubs #("Tracklet") VMS_L5D3PHI1Z1n1(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z1n1),
.enable(VMR_L5D3_VMS_L5D3PHI1Z1n1_wr_en),
.number_out(VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_number),
.read_add(VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_read_add),
.data_out(VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI1Z1n1;
wire VMR_L6D3_VMS_L6D3PHI1Z1n1_wr_en;
wire [5:0] VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_number;
wire [10:0] VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_read_add;
wire [17:0] VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1;
VMStubs #("Tracklet") VMS_L6D3PHI1Z1n1(
.data_in(VMR_L6D3_VMS_L6D3PHI1Z1n1),
.enable(VMR_L6D3_VMS_L6D3PHI1Z1n1_wr_en),
.number_out(VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_number),
.read_add(VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_read_add),
.data_out(VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z1n2;
wire VMR_L5D3_VMS_L5D3PHI1Z1n2_wr_en;
wire [5:0] VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1_number;
wire [10:0] VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1_read_add;
wire [17:0] VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1;
VMStubs #("Tracklet") VMS_L5D3PHI1Z1n2(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z1n2),
.enable(VMR_L5D3_VMS_L5D3PHI1Z1n2_wr_en),
.number_out(VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1_number),
.read_add(VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1_read_add),
.data_out(VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z1n1;
wire VMR_L6D3_VMS_L6D3PHI2Z1n1_wr_en;
wire [5:0] VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1_number;
wire [10:0] VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1_read_add;
wire [17:0] VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1;
VMStubs #("Tracklet") VMS_L6D3PHI2Z1n1(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z1n1),
.enable(VMR_L6D3_VMS_L6D3PHI2Z1n1_wr_en),
.number_out(VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1_number),
.read_add(VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1_read_add),
.data_out(VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z1n1;
wire VMR_L5D3_VMS_L5D3PHI2Z1n1_wr_en;
wire [5:0] VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1_number;
wire [10:0] VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1_read_add;
wire [17:0] VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1;
VMStubs #("Tracklet") VMS_L5D3PHI2Z1n1(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z1n1),
.enable(VMR_L5D3_VMS_L5D3PHI2Z1n1_wr_en),
.number_out(VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1_number),
.read_add(VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1_read_add),
.data_out(VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z1n2;
wire VMR_L6D3_VMS_L6D3PHI2Z1n2_wr_en;
wire [5:0] VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1_number;
wire [10:0] VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1_read_add;
wire [17:0] VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1;
VMStubs #("Tracklet") VMS_L6D3PHI2Z1n2(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z1n2),
.enable(VMR_L6D3_VMS_L6D3PHI2Z1n2_wr_en),
.number_out(VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1_number),
.read_add(VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1_read_add),
.data_out(VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z1n2;
wire VMR_L5D3_VMS_L5D3PHI2Z1n2_wr_en;
wire [5:0] VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1_number;
wire [10:0] VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1_read_add;
wire [17:0] VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1;
VMStubs #("Tracklet") VMS_L5D3PHI2Z1n2(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z1n2),
.enable(VMR_L5D3_VMS_L5D3PHI2Z1n2_wr_en),
.number_out(VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1_number),
.read_add(VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1_read_add),
.data_out(VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z1n1;
wire VMR_L6D3_VMS_L6D3PHI3Z1n1_wr_en;
wire [5:0] VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1_number;
wire [10:0] VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1_read_add;
wire [17:0] VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1;
VMStubs #("Tracklet") VMS_L6D3PHI3Z1n1(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z1n1),
.enable(VMR_L6D3_VMS_L6D3PHI3Z1n1_wr_en),
.number_out(VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1_number),
.read_add(VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1_read_add),
.data_out(VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z1n1;
wire VMR_L5D3_VMS_L5D3PHI3Z1n1_wr_en;
wire [5:0] VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1_number;
wire [10:0] VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1_read_add;
wire [17:0] VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1;
VMStubs #("Tracklet") VMS_L5D3PHI3Z1n1(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z1n1),
.enable(VMR_L5D3_VMS_L5D3PHI3Z1n1_wr_en),
.number_out(VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1_number),
.read_add(VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1_read_add),
.data_out(VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z1n2;
wire VMR_L6D3_VMS_L6D3PHI3Z1n2_wr_en;
wire [5:0] VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1_number;
wire [10:0] VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1_read_add;
wire [17:0] VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1;
VMStubs #("Tracklet") VMS_L6D3PHI3Z1n2(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z1n2),
.enable(VMR_L6D3_VMS_L6D3PHI3Z1n2_wr_en),
.number_out(VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1_number),
.read_add(VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1_read_add),
.data_out(VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z1n2;
wire VMR_L5D3_VMS_L5D3PHI3Z1n2_wr_en;
wire [5:0] VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1_number;
wire [10:0] VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1_read_add;
wire [17:0] VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1;
VMStubs #("Tracklet") VMS_L5D3PHI3Z1n2(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z1n2),
.enable(VMR_L5D3_VMS_L5D3PHI3Z1n2_wr_en),
.number_out(VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1_number),
.read_add(VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1_read_add),
.data_out(VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI4Z1n1;
wire VMR_L6D3_VMS_L6D3PHI4Z1n1_wr_en;
wire [5:0] VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1_number;
wire [10:0] VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1_read_add;
wire [17:0] VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1;
VMStubs #("Tracklet") VMS_L6D3PHI4Z1n1(
.data_in(VMR_L6D3_VMS_L6D3PHI4Z1n1),
.enable(VMR_L6D3_VMS_L6D3PHI4Z1n1_wr_en),
.number_out(VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1_number),
.read_add(VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1_read_add),
.data_out(VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z1n3;
wire VMR_L5D3_VMS_L5D3PHI1Z1n3_wr_en;
wire [5:0] VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2_number;
wire [10:0] VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2_read_add;
wire [17:0] VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2;
VMStubs #("Tracklet") VMS_L5D3PHI1Z1n3(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z1n3),
.enable(VMR_L5D3_VMS_L5D3PHI1Z1n3_wr_en),
.number_out(VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2_number),
.read_add(VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2_read_add),
.data_out(VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI1Z2n1;
wire VMR_L6D3_VMS_L6D3PHI1Z2n1_wr_en;
wire [5:0] VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2_number;
wire [10:0] VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2_read_add;
wire [17:0] VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2;
VMStubs #("Tracklet") VMS_L6D3PHI1Z2n1(
.data_in(VMR_L6D3_VMS_L6D3PHI1Z2n1),
.enable(VMR_L6D3_VMS_L6D3PHI1Z2n1_wr_en),
.number_out(VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2_number),
.read_add(VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2_read_add),
.data_out(VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z1n4;
wire VMR_L5D3_VMS_L5D3PHI1Z1n4_wr_en;
wire [5:0] VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2_number;
wire [10:0] VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2;
VMStubs #("Tracklet") VMS_L5D3PHI1Z1n4(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z1n4),
.enable(VMR_L5D3_VMS_L5D3PHI1Z1n4_wr_en),
.number_out(VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2_number),
.read_add(VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2_read_add),
.data_out(VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z2n1;
wire VMR_L6D3_VMS_L6D3PHI2Z2n1_wr_en;
wire [5:0] VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2_number;
wire [10:0] VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2;
VMStubs #("Tracklet") VMS_L6D3PHI2Z2n1(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z2n1),
.enable(VMR_L6D3_VMS_L6D3PHI2Z2n1_wr_en),
.number_out(VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2_number),
.read_add(VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2_read_add),
.data_out(VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z1n3;
wire VMR_L5D3_VMS_L5D3PHI2Z1n3_wr_en;
wire [5:0] VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2_number;
wire [10:0] VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2;
VMStubs #("Tracklet") VMS_L5D3PHI2Z1n3(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z1n3),
.enable(VMR_L5D3_VMS_L5D3PHI2Z1n3_wr_en),
.number_out(VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2_number),
.read_add(VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2_read_add),
.data_out(VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z2n2;
wire VMR_L6D3_VMS_L6D3PHI2Z2n2_wr_en;
wire [5:0] VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2_number;
wire [10:0] VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2;
VMStubs #("Tracklet") VMS_L6D3PHI2Z2n2(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z2n2),
.enable(VMR_L6D3_VMS_L6D3PHI2Z2n2_wr_en),
.number_out(VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2_number),
.read_add(VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2_read_add),
.data_out(VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z1n4;
wire VMR_L5D3_VMS_L5D3PHI2Z1n4_wr_en;
wire [5:0] VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2_number;
wire [10:0] VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2;
VMStubs #("Tracklet") VMS_L5D3PHI2Z1n4(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z1n4),
.enable(VMR_L5D3_VMS_L5D3PHI2Z1n4_wr_en),
.number_out(VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2_number),
.read_add(VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2_read_add),
.data_out(VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z2n1;
wire VMR_L6D3_VMS_L6D3PHI3Z2n1_wr_en;
wire [5:0] VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2_number;
wire [10:0] VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2;
VMStubs #("Tracklet") VMS_L6D3PHI3Z2n1(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z2n1),
.enable(VMR_L6D3_VMS_L6D3PHI3Z2n1_wr_en),
.number_out(VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2_number),
.read_add(VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2_read_add),
.data_out(VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z1n3;
wire VMR_L5D3_VMS_L5D3PHI3Z1n3_wr_en;
wire [5:0] VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2_number;
wire [10:0] VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2;
VMStubs #("Tracklet") VMS_L5D3PHI3Z1n3(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z1n3),
.enable(VMR_L5D3_VMS_L5D3PHI3Z1n3_wr_en),
.number_out(VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2_number),
.read_add(VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2_read_add),
.data_out(VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z2n2;
wire VMR_L6D3_VMS_L6D3PHI3Z2n2_wr_en;
wire [5:0] VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2_number;
wire [10:0] VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2;
VMStubs #("Tracklet") VMS_L6D3PHI3Z2n2(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z2n2),
.enable(VMR_L6D3_VMS_L6D3PHI3Z2n2_wr_en),
.number_out(VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2_number),
.read_add(VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2_read_add),
.data_out(VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z1n4;
wire VMR_L5D3_VMS_L5D3PHI3Z1n4_wr_en;
wire [5:0] VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2_number;
wire [10:0] VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2_read_add;
wire [17:0] VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2;
VMStubs #("Tracklet") VMS_L5D3PHI3Z1n4(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z1n4),
.enable(VMR_L5D3_VMS_L5D3PHI3Z1n4_wr_en),
.number_out(VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2_number),
.read_add(VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2_read_add),
.data_out(VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI4Z2n1;
wire VMR_L6D3_VMS_L6D3PHI4Z2n1_wr_en;
wire [5:0] VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2_number;
wire [10:0] VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2_read_add;
wire [17:0] VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2;
VMStubs #("Tracklet") VMS_L6D3PHI4Z2n1(
.data_in(VMR_L6D3_VMS_L6D3PHI4Z2n1),
.enable(VMR_L6D3_VMS_L6D3PHI4Z2n1_wr_en),
.number_out(VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2_number),
.read_add(VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2_read_add),
.data_out(VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z2n1;
wire VMR_L5D3_VMS_L5D3PHI1Z2n1_wr_en;
wire [5:0] VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2_number;
wire [10:0] VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2_read_add;
wire [17:0] VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2;
VMStubs #("Tracklet") VMS_L5D3PHI1Z2n1(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z2n1),
.enable(VMR_L5D3_VMS_L5D3PHI1Z2n1_wr_en),
.number_out(VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2_number),
.read_add(VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2_read_add),
.data_out(VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI1Z2n2;
wire VMR_L6D3_VMS_L6D3PHI1Z2n2_wr_en;
wire [5:0] VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2_number;
wire [10:0] VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2_read_add;
wire [17:0] VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2;
VMStubs #("Tracklet") VMS_L6D3PHI1Z2n2(
.data_in(VMR_L6D3_VMS_L6D3PHI1Z2n2),
.enable(VMR_L6D3_VMS_L6D3PHI1Z2n2_wr_en),
.number_out(VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2_number),
.read_add(VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2_read_add),
.data_out(VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z2n2;
wire VMR_L5D3_VMS_L5D3PHI1Z2n2_wr_en;
wire [5:0] VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2_number;
wire [10:0] VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2;
VMStubs #("Tracklet") VMS_L5D3PHI1Z2n2(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z2n2),
.enable(VMR_L5D3_VMS_L5D3PHI1Z2n2_wr_en),
.number_out(VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2_number),
.read_add(VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2_read_add),
.data_out(VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z2n3;
wire VMR_L6D3_VMS_L6D3PHI2Z2n3_wr_en;
wire [5:0] VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2_number;
wire [10:0] VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2;
VMStubs #("Tracklet") VMS_L6D3PHI2Z2n3(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z2n3),
.enable(VMR_L6D3_VMS_L6D3PHI2Z2n3_wr_en),
.number_out(VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2_number),
.read_add(VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2_read_add),
.data_out(VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z2n1;
wire VMR_L5D3_VMS_L5D3PHI2Z2n1_wr_en;
wire [5:0] VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2_number;
wire [10:0] VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2;
VMStubs #("Tracklet") VMS_L5D3PHI2Z2n1(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z2n1),
.enable(VMR_L5D3_VMS_L5D3PHI2Z2n1_wr_en),
.number_out(VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2_number),
.read_add(VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2_read_add),
.data_out(VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z2n4;
wire VMR_L6D3_VMS_L6D3PHI2Z2n4_wr_en;
wire [5:0] VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2_number;
wire [10:0] VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2;
VMStubs #("Tracklet") VMS_L6D3PHI2Z2n4(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z2n4),
.enable(VMR_L6D3_VMS_L6D3PHI2Z2n4_wr_en),
.number_out(VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2_number),
.read_add(VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2_read_add),
.data_out(VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z2n2;
wire VMR_L5D3_VMS_L5D3PHI2Z2n2_wr_en;
wire [5:0] VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2_number;
wire [10:0] VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2;
VMStubs #("Tracklet") VMS_L5D3PHI2Z2n2(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z2n2),
.enable(VMR_L5D3_VMS_L5D3PHI2Z2n2_wr_en),
.number_out(VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2_number),
.read_add(VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2_read_add),
.data_out(VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z2n3;
wire VMR_L6D3_VMS_L6D3PHI3Z2n3_wr_en;
wire [5:0] VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2_number;
wire [10:0] VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2;
VMStubs #("Tracklet") VMS_L6D3PHI3Z2n3(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z2n3),
.enable(VMR_L6D3_VMS_L6D3PHI3Z2n3_wr_en),
.number_out(VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2_number),
.read_add(VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2_read_add),
.data_out(VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z2n1;
wire VMR_L5D3_VMS_L5D3PHI3Z2n1_wr_en;
wire [5:0] VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2_number;
wire [10:0] VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2;
VMStubs #("Tracklet") VMS_L5D3PHI3Z2n1(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z2n1),
.enable(VMR_L5D3_VMS_L5D3PHI3Z2n1_wr_en),
.number_out(VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2_number),
.read_add(VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2_read_add),
.data_out(VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z2n4;
wire VMR_L6D3_VMS_L6D3PHI3Z2n4_wr_en;
wire [5:0] VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2_number;
wire [10:0] VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2;
VMStubs #("Tracklet") VMS_L6D3PHI3Z2n4(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z2n4),
.enable(VMR_L6D3_VMS_L6D3PHI3Z2n4_wr_en),
.number_out(VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2_number),
.read_add(VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2_read_add),
.data_out(VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z2n2;
wire VMR_L5D3_VMS_L5D3PHI3Z2n2_wr_en;
wire [5:0] VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_number;
wire [10:0] VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_read_add;
wire [17:0] VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2;
VMStubs #("Tracklet") VMS_L5D3PHI3Z2n2(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z2n2),
.enable(VMR_L5D3_VMS_L5D3PHI3Z2n2_wr_en),
.number_out(VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_number),
.read_add(VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_read_add),
.data_out(VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI4Z2n2;
wire VMR_L6D3_VMS_L6D3PHI4Z2n2_wr_en;
wire [5:0] VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_number;
wire [10:0] VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_read_add;
wire [17:0] VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2;
VMStubs #("Tracklet") VMS_L6D3PHI4Z2n2(
.data_in(VMR_L6D3_VMS_L6D3PHI4Z2n2),
.enable(VMR_L6D3_VMS_L6D3PHI4Z2n2_wr_en),
.number_out(VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_number),
.read_add(VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_read_add),
.data_out(VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z2n3;
wire VMR_L5D3_VMS_L5D3PHI1Z2n3_wr_en;
wire [5:0] VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1_number;
wire [10:0] VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1_read_add;
wire [17:0] VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1;
VMStubs #("Tracklet") VMS_L5D3PHI1Z2n3(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z2n3),
.enable(VMR_L5D3_VMS_L5D3PHI1Z2n3_wr_en),
.number_out(VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1_number),
.read_add(VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1_read_add),
.data_out(VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI1Z1n1;
wire VMR_L6D4_VMS_L6D4PHI1Z1n1_wr_en;
wire [5:0] VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1_number;
wire [10:0] VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1_read_add;
wire [17:0] VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1;
VMStubs #("Tracklet") VMS_L6D4PHI1Z1n1(
.data_in(VMR_L6D4_VMS_L6D4PHI1Z1n1),
.enable(VMR_L6D4_VMS_L6D4PHI1Z1n1_wr_en),
.number_out(VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1_number),
.read_add(VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1_read_add),
.data_out(VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z2n4;
wire VMR_L5D3_VMS_L5D3PHI1Z2n4_wr_en;
wire [5:0] VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1_number;
wire [10:0] VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1;
VMStubs #("Tracklet") VMS_L5D3PHI1Z2n4(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z2n4),
.enable(VMR_L5D3_VMS_L5D3PHI1Z2n4_wr_en),
.number_out(VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1_number),
.read_add(VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1_read_add),
.data_out(VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z1n1;
wire VMR_L6D4_VMS_L6D4PHI2Z1n1_wr_en;
wire [5:0] VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1_number;
wire [10:0] VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1;
VMStubs #("Tracklet") VMS_L6D4PHI2Z1n1(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z1n1),
.enable(VMR_L6D4_VMS_L6D4PHI2Z1n1_wr_en),
.number_out(VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1_number),
.read_add(VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1_read_add),
.data_out(VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z2n3;
wire VMR_L5D3_VMS_L5D3PHI2Z2n3_wr_en;
wire [5:0] VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1_number;
wire [10:0] VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1;
VMStubs #("Tracklet") VMS_L5D3PHI2Z2n3(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z2n3),
.enable(VMR_L5D3_VMS_L5D3PHI2Z2n3_wr_en),
.number_out(VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1_number),
.read_add(VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1_read_add),
.data_out(VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z1n2;
wire VMR_L6D4_VMS_L6D4PHI2Z1n2_wr_en;
wire [5:0] VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1_number;
wire [10:0] VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1;
VMStubs #("Tracklet") VMS_L6D4PHI2Z1n2(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z1n2),
.enable(VMR_L6D4_VMS_L6D4PHI2Z1n2_wr_en),
.number_out(VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1_number),
.read_add(VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1_read_add),
.data_out(VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z2n4;
wire VMR_L5D3_VMS_L5D3PHI2Z2n4_wr_en;
wire [5:0] VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1_number;
wire [10:0] VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1;
VMStubs #("Tracklet") VMS_L5D3PHI2Z2n4(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z2n4),
.enable(VMR_L5D3_VMS_L5D3PHI2Z2n4_wr_en),
.number_out(VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1_number),
.read_add(VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1_read_add),
.data_out(VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z1n1;
wire VMR_L6D4_VMS_L6D4PHI3Z1n1_wr_en;
wire [5:0] VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1_number;
wire [10:0] VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1;
VMStubs #("Tracklet") VMS_L6D4PHI3Z1n1(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z1n1),
.enable(VMR_L6D4_VMS_L6D4PHI3Z1n1_wr_en),
.number_out(VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1_number),
.read_add(VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1_read_add),
.data_out(VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z2n3;
wire VMR_L5D3_VMS_L5D3PHI3Z2n3_wr_en;
wire [5:0] VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1_number;
wire [10:0] VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1;
VMStubs #("Tracklet") VMS_L5D3PHI3Z2n3(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z2n3),
.enable(VMR_L5D3_VMS_L5D3PHI3Z2n3_wr_en),
.number_out(VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1_number),
.read_add(VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1_read_add),
.data_out(VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z1n2;
wire VMR_L6D4_VMS_L6D4PHI3Z1n2_wr_en;
wire [5:0] VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1_number;
wire [10:0] VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1;
VMStubs #("Tracklet") VMS_L6D4PHI3Z1n2(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z1n2),
.enable(VMR_L6D4_VMS_L6D4PHI3Z1n2_wr_en),
.number_out(VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1_number),
.read_add(VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1_read_add),
.data_out(VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z2n4;
wire VMR_L5D3_VMS_L5D3PHI3Z2n4_wr_en;
wire [5:0] VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1_number;
wire [10:0] VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1_read_add;
wire [17:0] VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1;
VMStubs #("Tracklet") VMS_L5D3PHI3Z2n4(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z2n4),
.enable(VMR_L5D3_VMS_L5D3PHI3Z2n4_wr_en),
.number_out(VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1_number),
.read_add(VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1_read_add),
.data_out(VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI4Z1n1;
wire VMR_L6D4_VMS_L6D4PHI4Z1n1_wr_en;
wire [5:0] VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1_number;
wire [10:0] VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1_read_add;
wire [17:0] VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1;
VMStubs #("Tracklet") VMS_L6D4PHI4Z1n1(
.data_in(VMR_L6D4_VMS_L6D4PHI4Z1n1),
.enable(VMR_L6D4_VMS_L6D4PHI4Z1n1_wr_en),
.number_out(VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1_number),
.read_add(VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1_read_add),
.data_out(VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z1n1;
wire VMR_L5D4_VMS_L5D4PHI1Z1n1_wr_en;
wire [5:0] VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1_number;
wire [10:0] VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1_read_add;
wire [17:0] VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1;
VMStubs #("Tracklet") VMS_L5D4PHI1Z1n1(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z1n1),
.enable(VMR_L5D4_VMS_L5D4PHI1Z1n1_wr_en),
.number_out(VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1_number),
.read_add(VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1_read_add),
.data_out(VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI1Z1n2;
wire VMR_L6D4_VMS_L6D4PHI1Z1n2_wr_en;
wire [5:0] VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1_number;
wire [10:0] VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1_read_add;
wire [17:0] VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1;
VMStubs #("Tracklet") VMS_L6D4PHI1Z1n2(
.data_in(VMR_L6D4_VMS_L6D4PHI1Z1n2),
.enable(VMR_L6D4_VMS_L6D4PHI1Z1n2_wr_en),
.number_out(VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1_number),
.read_add(VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1_read_add),
.data_out(VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z1n2;
wire VMR_L5D4_VMS_L5D4PHI1Z1n2_wr_en;
wire [5:0] VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1_number;
wire [10:0] VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1;
VMStubs #("Tracklet") VMS_L5D4PHI1Z1n2(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z1n2),
.enable(VMR_L5D4_VMS_L5D4PHI1Z1n2_wr_en),
.number_out(VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1_number),
.read_add(VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1_read_add),
.data_out(VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z1n3;
wire VMR_L6D4_VMS_L6D4PHI2Z1n3_wr_en;
wire [5:0] VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1_number;
wire [10:0] VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1;
VMStubs #("Tracklet") VMS_L6D4PHI2Z1n3(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z1n3),
.enable(VMR_L6D4_VMS_L6D4PHI2Z1n3_wr_en),
.number_out(VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1_number),
.read_add(VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1_read_add),
.data_out(VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z1n1;
wire VMR_L5D4_VMS_L5D4PHI2Z1n1_wr_en;
wire [5:0] VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1_number;
wire [10:0] VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1;
VMStubs #("Tracklet") VMS_L5D4PHI2Z1n1(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z1n1),
.enable(VMR_L5D4_VMS_L5D4PHI2Z1n1_wr_en),
.number_out(VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1_number),
.read_add(VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1_read_add),
.data_out(VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z1n4;
wire VMR_L6D4_VMS_L6D4PHI2Z1n4_wr_en;
wire [5:0] VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1_number;
wire [10:0] VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1;
VMStubs #("Tracklet") VMS_L6D4PHI2Z1n4(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z1n4),
.enable(VMR_L6D4_VMS_L6D4PHI2Z1n4_wr_en),
.number_out(VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1_number),
.read_add(VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1_read_add),
.data_out(VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z1n2;
wire VMR_L5D4_VMS_L5D4PHI2Z1n2_wr_en;
wire [5:0] VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1_number;
wire [10:0] VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1;
VMStubs #("Tracklet") VMS_L5D4PHI2Z1n2(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z1n2),
.enable(VMR_L5D4_VMS_L5D4PHI2Z1n2_wr_en),
.number_out(VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1_number),
.read_add(VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1_read_add),
.data_out(VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z1n3;
wire VMR_L6D4_VMS_L6D4PHI3Z1n3_wr_en;
wire [5:0] VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1_number;
wire [10:0] VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1;
VMStubs #("Tracklet") VMS_L6D4PHI3Z1n3(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z1n3),
.enable(VMR_L6D4_VMS_L6D4PHI3Z1n3_wr_en),
.number_out(VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1_number),
.read_add(VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1_read_add),
.data_out(VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z1n1;
wire VMR_L5D4_VMS_L5D4PHI3Z1n1_wr_en;
wire [5:0] VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1_number;
wire [10:0] VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1;
VMStubs #("Tracklet") VMS_L5D4PHI3Z1n1(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z1n1),
.enable(VMR_L5D4_VMS_L5D4PHI3Z1n1_wr_en),
.number_out(VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1_number),
.read_add(VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1_read_add),
.data_out(VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z1n4;
wire VMR_L6D4_VMS_L6D4PHI3Z1n4_wr_en;
wire [5:0] VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1_number;
wire [10:0] VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1;
VMStubs #("Tracklet") VMS_L6D4PHI3Z1n4(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z1n4),
.enable(VMR_L6D4_VMS_L6D4PHI3Z1n4_wr_en),
.number_out(VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1_number),
.read_add(VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1_read_add),
.data_out(VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z1n2;
wire VMR_L5D4_VMS_L5D4PHI3Z1n2_wr_en;
wire [5:0] VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_number;
wire [10:0] VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_read_add;
wire [17:0] VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1;
VMStubs #("Tracklet") VMS_L5D4PHI3Z1n2(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z1n2),
.enable(VMR_L5D4_VMS_L5D4PHI3Z1n2_wr_en),
.number_out(VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_number),
.read_add(VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_read_add),
.data_out(VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI4Z1n2;
wire VMR_L6D4_VMS_L6D4PHI4Z1n2_wr_en;
wire [5:0] VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_number;
wire [10:0] VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_read_add;
wire [17:0] VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1;
VMStubs #("Tracklet") VMS_L6D4PHI4Z1n2(
.data_in(VMR_L6D4_VMS_L6D4PHI4Z1n2),
.enable(VMR_L6D4_VMS_L6D4PHI4Z1n2_wr_en),
.number_out(VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_number),
.read_add(VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_read_add),
.data_out(VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z1n3;
wire VMR_L5D4_VMS_L5D4PHI1Z1n3_wr_en;
wire [5:0] VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2_number;
wire [10:0] VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2_read_add;
wire [17:0] VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2;
VMStubs #("Tracklet") VMS_L5D4PHI1Z1n3(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z1n3),
.enable(VMR_L5D4_VMS_L5D4PHI1Z1n3_wr_en),
.number_out(VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2_number),
.read_add(VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2_read_add),
.data_out(VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI1Z2n1;
wire VMR_L6D4_VMS_L6D4PHI1Z2n1_wr_en;
wire [5:0] VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2_number;
wire [10:0] VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2_read_add;
wire [17:0] VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2;
VMStubs #("Tracklet") VMS_L6D4PHI1Z2n1(
.data_in(VMR_L6D4_VMS_L6D4PHI1Z2n1),
.enable(VMR_L6D4_VMS_L6D4PHI1Z2n1_wr_en),
.number_out(VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2_number),
.read_add(VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2_read_add),
.data_out(VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z1n4;
wire VMR_L5D4_VMS_L5D4PHI1Z1n4_wr_en;
wire [5:0] VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2_number;
wire [10:0] VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2;
VMStubs #("Tracklet") VMS_L5D4PHI1Z1n4(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z1n4),
.enable(VMR_L5D4_VMS_L5D4PHI1Z1n4_wr_en),
.number_out(VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2_number),
.read_add(VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2_read_add),
.data_out(VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z2n1;
wire VMR_L6D4_VMS_L6D4PHI2Z2n1_wr_en;
wire [5:0] VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2_number;
wire [10:0] VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2;
VMStubs #("Tracklet") VMS_L6D4PHI2Z2n1(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z2n1),
.enable(VMR_L6D4_VMS_L6D4PHI2Z2n1_wr_en),
.number_out(VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2_number),
.read_add(VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2_read_add),
.data_out(VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z1n3;
wire VMR_L5D4_VMS_L5D4PHI2Z1n3_wr_en;
wire [5:0] VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2_number;
wire [10:0] VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2;
VMStubs #("Tracklet") VMS_L5D4PHI2Z1n3(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z1n3),
.enable(VMR_L5D4_VMS_L5D4PHI2Z1n3_wr_en),
.number_out(VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2_number),
.read_add(VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2_read_add),
.data_out(VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z2n2;
wire VMR_L6D4_VMS_L6D4PHI2Z2n2_wr_en;
wire [5:0] VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2_number;
wire [10:0] VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2;
VMStubs #("Tracklet") VMS_L6D4PHI2Z2n2(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z2n2),
.enable(VMR_L6D4_VMS_L6D4PHI2Z2n2_wr_en),
.number_out(VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2_number),
.read_add(VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2_read_add),
.data_out(VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z1n4;
wire VMR_L5D4_VMS_L5D4PHI2Z1n4_wr_en;
wire [5:0] VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2_number;
wire [10:0] VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2;
VMStubs #("Tracklet") VMS_L5D4PHI2Z1n4(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z1n4),
.enable(VMR_L5D4_VMS_L5D4PHI2Z1n4_wr_en),
.number_out(VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2_number),
.read_add(VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2_read_add),
.data_out(VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z2n1;
wire VMR_L6D4_VMS_L6D4PHI3Z2n1_wr_en;
wire [5:0] VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2_number;
wire [10:0] VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2;
VMStubs #("Tracklet") VMS_L6D4PHI3Z2n1(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z2n1),
.enable(VMR_L6D4_VMS_L6D4PHI3Z2n1_wr_en),
.number_out(VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2_number),
.read_add(VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2_read_add),
.data_out(VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z1n3;
wire VMR_L5D4_VMS_L5D4PHI3Z1n3_wr_en;
wire [5:0] VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2_number;
wire [10:0] VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2;
VMStubs #("Tracklet") VMS_L5D4PHI3Z1n3(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z1n3),
.enable(VMR_L5D4_VMS_L5D4PHI3Z1n3_wr_en),
.number_out(VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2_number),
.read_add(VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2_read_add),
.data_out(VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z2n2;
wire VMR_L6D4_VMS_L6D4PHI3Z2n2_wr_en;
wire [5:0] VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2_number;
wire [10:0] VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2;
VMStubs #("Tracklet") VMS_L6D4PHI3Z2n2(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z2n2),
.enable(VMR_L6D4_VMS_L6D4PHI3Z2n2_wr_en),
.number_out(VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2_number),
.read_add(VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2_read_add),
.data_out(VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z1n4;
wire VMR_L5D4_VMS_L5D4PHI3Z1n4_wr_en;
wire [5:0] VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2_number;
wire [10:0] VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2_read_add;
wire [17:0] VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2;
VMStubs #("Tracklet") VMS_L5D4PHI3Z1n4(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z1n4),
.enable(VMR_L5D4_VMS_L5D4PHI3Z1n4_wr_en),
.number_out(VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2_number),
.read_add(VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2_read_add),
.data_out(VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI4Z2n1;
wire VMR_L6D4_VMS_L6D4PHI4Z2n1_wr_en;
wire [5:0] VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2_number;
wire [10:0] VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2_read_add;
wire [17:0] VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2;
VMStubs #("Tracklet") VMS_L6D4PHI4Z2n1(
.data_in(VMR_L6D4_VMS_L6D4PHI4Z2n1),
.enable(VMR_L6D4_VMS_L6D4PHI4Z2n1_wr_en),
.number_out(VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2_number),
.read_add(VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2_read_add),
.data_out(VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z2n1;
wire VMR_L5D4_VMS_L5D4PHI1Z2n1_wr_en;
wire [5:0] VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2_number;
wire [10:0] VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2_read_add;
wire [17:0] VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2;
VMStubs #("Tracklet") VMS_L5D4PHI1Z2n1(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z2n1),
.enable(VMR_L5D4_VMS_L5D4PHI1Z2n1_wr_en),
.number_out(VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2_number),
.read_add(VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2_read_add),
.data_out(VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI1Z2n2;
wire VMR_L6D4_VMS_L6D4PHI1Z2n2_wr_en;
wire [5:0] VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2_number;
wire [10:0] VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2_read_add;
wire [17:0] VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2;
VMStubs #("Tracklet") VMS_L6D4PHI1Z2n2(
.data_in(VMR_L6D4_VMS_L6D4PHI1Z2n2),
.enable(VMR_L6D4_VMS_L6D4PHI1Z2n2_wr_en),
.number_out(VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2_number),
.read_add(VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2_read_add),
.data_out(VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z2n2;
wire VMR_L5D4_VMS_L5D4PHI1Z2n2_wr_en;
wire [5:0] VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2_number;
wire [10:0] VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2;
VMStubs #("Tracklet") VMS_L5D4PHI1Z2n2(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z2n2),
.enable(VMR_L5D4_VMS_L5D4PHI1Z2n2_wr_en),
.number_out(VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2_number),
.read_add(VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2_read_add),
.data_out(VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z2n3;
wire VMR_L6D4_VMS_L6D4PHI2Z2n3_wr_en;
wire [5:0] VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2_number;
wire [10:0] VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2;
VMStubs #("Tracklet") VMS_L6D4PHI2Z2n3(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z2n3),
.enable(VMR_L6D4_VMS_L6D4PHI2Z2n3_wr_en),
.number_out(VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2_number),
.read_add(VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2_read_add),
.data_out(VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z2n1;
wire VMR_L5D4_VMS_L5D4PHI2Z2n1_wr_en;
wire [5:0] VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2_number;
wire [10:0] VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2;
VMStubs #("Tracklet") VMS_L5D4PHI2Z2n1(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z2n1),
.enable(VMR_L5D4_VMS_L5D4PHI2Z2n1_wr_en),
.number_out(VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2_number),
.read_add(VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2_read_add),
.data_out(VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z2n4;
wire VMR_L6D4_VMS_L6D4PHI2Z2n4_wr_en;
wire [5:0] VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2_number;
wire [10:0] VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2;
VMStubs #("Tracklet") VMS_L6D4PHI2Z2n4(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z2n4),
.enable(VMR_L6D4_VMS_L6D4PHI2Z2n4_wr_en),
.number_out(VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2_number),
.read_add(VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2_read_add),
.data_out(VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z2n2;
wire VMR_L5D4_VMS_L5D4PHI2Z2n2_wr_en;
wire [5:0] VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2_number;
wire [10:0] VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2;
VMStubs #("Tracklet") VMS_L5D4PHI2Z2n2(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z2n2),
.enable(VMR_L5D4_VMS_L5D4PHI2Z2n2_wr_en),
.number_out(VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2_number),
.read_add(VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2_read_add),
.data_out(VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z2n3;
wire VMR_L6D4_VMS_L6D4PHI3Z2n3_wr_en;
wire [5:0] VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2_number;
wire [10:0] VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2;
VMStubs #("Tracklet") VMS_L6D4PHI3Z2n3(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z2n3),
.enable(VMR_L6D4_VMS_L6D4PHI3Z2n3_wr_en),
.number_out(VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2_number),
.read_add(VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2_read_add),
.data_out(VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z2n1;
wire VMR_L5D4_VMS_L5D4PHI3Z2n1_wr_en;
wire [5:0] VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2_number;
wire [10:0] VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2;
VMStubs #("Tracklet") VMS_L5D4PHI3Z2n1(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z2n1),
.enable(VMR_L5D4_VMS_L5D4PHI3Z2n1_wr_en),
.number_out(VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2_number),
.read_add(VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2_read_add),
.data_out(VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z2n4;
wire VMR_L6D4_VMS_L6D4PHI3Z2n4_wr_en;
wire [5:0] VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2_number;
wire [10:0] VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2;
VMStubs #("Tracklet") VMS_L6D4PHI3Z2n4(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z2n4),
.enable(VMR_L6D4_VMS_L6D4PHI3Z2n4_wr_en),
.number_out(VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2_number),
.read_add(VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2_read_add),
.data_out(VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z2n2;
wire VMR_L5D4_VMS_L5D4PHI3Z2n2_wr_en;
wire [5:0] VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_number;
wire [10:0] VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_read_add;
wire [17:0] VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2;
VMStubs #("Tracklet") VMS_L5D4PHI3Z2n2(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z2n2),
.enable(VMR_L5D4_VMS_L5D4PHI3Z2n2_wr_en),
.number_out(VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_number),
.read_add(VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_read_add),
.data_out(VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI4Z2n2;
wire VMR_L6D4_VMS_L6D4PHI4Z2n2_wr_en;
wire [5:0] VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_number;
wire [10:0] VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_read_add;
wire [17:0] VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2;
VMStubs #("Tracklet") VMS_L6D4PHI4Z2n2(
.data_in(VMR_L6D4_VMS_L6D4PHI4Z2n2),
.enable(VMR_L6D4_VMS_L6D4PHI4Z2n2_wr_en),
.number_out(VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_number),
.read_add(VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_read_add),
.data_out(VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z1_L2D3PHI1Z1_SP_L1D3PHI1Z1_L2D3PHI1Z1;
wire TE_L1D3PHI1Z1_L2D3PHI1Z1_SP_L1D3PHI1Z1_L2D3PHI1Z1_wr_en;
wire [5:0] SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1Z1_L2D3PHI1Z1(
.data_in(TE_L1D3PHI1Z1_L2D3PHI1Z1_SP_L1D3PHI1Z1_L2D3PHI1Z1),
.enable(TE_L1D3PHI1Z1_L2D3PHI1Z1_SP_L1D3PHI1Z1_L2D3PHI1Z1_wr_en),
.number_out(SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3),
.start(start4_0),
.done(done3_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z1_L2D3PHI2Z1_SP_L1D3PHI1Z1_L2D3PHI2Z1;
wire TE_L1D3PHI1Z1_L2D3PHI2Z1_SP_L1D3PHI1Z1_L2D3PHI2Z1_wr_en;
wire [5:0] SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1Z1_L2D3PHI2Z1(
.data_in(TE_L1D3PHI1Z1_L2D3PHI2Z1_SP_L1D3PHI1Z1_L2D3PHI2Z1),
.enable(TE_L1D3PHI1Z1_L2D3PHI2Z1_SP_L1D3PHI1Z1_L2D3PHI2Z1_wr_en),
.number_out(SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z1_L2D3PHI2Z1_SP_L1D3PHI2Z1_L2D3PHI2Z1;
wire TE_L1D3PHI2Z1_L2D3PHI2Z1_SP_L1D3PHI2Z1_L2D3PHI2Z1_wr_en;
wire [5:0] SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2Z1_L2D3PHI2Z1(
.data_in(TE_L1D3PHI2Z1_L2D3PHI2Z1_SP_L1D3PHI2Z1_L2D3PHI2Z1),
.enable(TE_L1D3PHI2Z1_L2D3PHI2Z1_SP_L1D3PHI2Z1_L2D3PHI2Z1_wr_en),
.number_out(SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z1_L2D3PHI3Z1_SP_L1D3PHI2Z1_L2D3PHI3Z1;
wire TE_L1D3PHI2Z1_L2D3PHI3Z1_SP_L1D3PHI2Z1_L2D3PHI3Z1_wr_en;
wire [5:0] SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2Z1_L2D3PHI3Z1(
.data_in(TE_L1D3PHI2Z1_L2D3PHI3Z1_SP_L1D3PHI2Z1_L2D3PHI3Z1),
.enable(TE_L1D3PHI2Z1_L2D3PHI3Z1_SP_L1D3PHI2Z1_L2D3PHI3Z1_wr_en),
.number_out(SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z1_L2D3PHI3Z1_SP_L1D3PHI3Z1_L2D3PHI3Z1;
wire TE_L1D3PHI3Z1_L2D3PHI3Z1_SP_L1D3PHI3Z1_L2D3PHI3Z1_wr_en;
wire [5:0] SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3Z1_L2D3PHI3Z1(
.data_in(TE_L1D3PHI3Z1_L2D3PHI3Z1_SP_L1D3PHI3Z1_L2D3PHI3Z1),
.enable(TE_L1D3PHI3Z1_L2D3PHI3Z1_SP_L1D3PHI3Z1_L2D3PHI3Z1_wr_en),
.number_out(SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z1_L2D3PHI4Z1_SP_L1D3PHI3Z1_L2D3PHI4Z1;
wire TE_L1D3PHI3Z1_L2D3PHI4Z1_SP_L1D3PHI3Z1_L2D3PHI4Z1_wr_en;
wire [5:0] SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3Z1_L2D3PHI4Z1(
.data_in(TE_L1D3PHI3Z1_L2D3PHI4Z1_SP_L1D3PHI3Z1_L2D3PHI4Z1),
.enable(TE_L1D3PHI3Z1_L2D3PHI4Z1_SP_L1D3PHI3Z1_L2D3PHI4Z1_wr_en),
.number_out(SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z1_L2D3PHI1Z2_SP_L1D3PHI1Z1_L2D3PHI1Z2;
wire TE_L1D3PHI1Z1_L2D3PHI1Z2_SP_L1D3PHI1Z1_L2D3PHI1Z2_wr_en;
wire [5:0] SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1Z1_L2D3PHI1Z2(
.data_in(TE_L1D3PHI1Z1_L2D3PHI1Z2_SP_L1D3PHI1Z1_L2D3PHI1Z2),
.enable(TE_L1D3PHI1Z1_L2D3PHI1Z2_SP_L1D3PHI1Z1_L2D3PHI1Z2_wr_en),
.number_out(SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z1_L2D3PHI2Z2_SP_L1D3PHI1Z1_L2D3PHI2Z2;
wire TE_L1D3PHI1Z1_L2D3PHI2Z2_SP_L1D3PHI1Z1_L2D3PHI2Z2_wr_en;
wire [5:0] SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1Z1_L2D3PHI2Z2(
.data_in(TE_L1D3PHI1Z1_L2D3PHI2Z2_SP_L1D3PHI1Z1_L2D3PHI2Z2),
.enable(TE_L1D3PHI1Z1_L2D3PHI2Z2_SP_L1D3PHI1Z1_L2D3PHI2Z2_wr_en),
.number_out(SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z1_L2D3PHI2Z2_SP_L1D3PHI2Z1_L2D3PHI2Z2;
wire TE_L1D3PHI2Z1_L2D3PHI2Z2_SP_L1D3PHI2Z1_L2D3PHI2Z2_wr_en;
wire [5:0] SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2Z1_L2D3PHI2Z2(
.data_in(TE_L1D3PHI2Z1_L2D3PHI2Z2_SP_L1D3PHI2Z1_L2D3PHI2Z2),
.enable(TE_L1D3PHI2Z1_L2D3PHI2Z2_SP_L1D3PHI2Z1_L2D3PHI2Z2_wr_en),
.number_out(SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z1_L2D3PHI3Z2_SP_L1D3PHI2Z1_L2D3PHI3Z2;
wire TE_L1D3PHI2Z1_L2D3PHI3Z2_SP_L1D3PHI2Z1_L2D3PHI3Z2_wr_en;
wire [5:0] SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2Z1_L2D3PHI3Z2(
.data_in(TE_L1D3PHI2Z1_L2D3PHI3Z2_SP_L1D3PHI2Z1_L2D3PHI3Z2),
.enable(TE_L1D3PHI2Z1_L2D3PHI3Z2_SP_L1D3PHI2Z1_L2D3PHI3Z2_wr_en),
.number_out(SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z1_L2D3PHI3Z2_SP_L1D3PHI3Z1_L2D3PHI3Z2;
wire TE_L1D3PHI3Z1_L2D3PHI3Z2_SP_L1D3PHI3Z1_L2D3PHI3Z2_wr_en;
wire [5:0] SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3Z1_L2D3PHI3Z2(
.data_in(TE_L1D3PHI3Z1_L2D3PHI3Z2_SP_L1D3PHI3Z1_L2D3PHI3Z2),
.enable(TE_L1D3PHI3Z1_L2D3PHI3Z2_SP_L1D3PHI3Z1_L2D3PHI3Z2_wr_en),
.number_out(SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z1_L2D3PHI4Z2_SP_L1D3PHI3Z1_L2D3PHI4Z2;
wire TE_L1D3PHI3Z1_L2D3PHI4Z2_SP_L1D3PHI3Z1_L2D3PHI4Z2_wr_en;
wire [5:0] SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3Z1_L2D3PHI4Z2(
.data_in(TE_L1D3PHI3Z1_L2D3PHI4Z2_SP_L1D3PHI3Z1_L2D3PHI4Z2),
.enable(TE_L1D3PHI3Z1_L2D3PHI4Z2_SP_L1D3PHI3Z1_L2D3PHI4Z2_wr_en),
.number_out(SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z2_L2D3PHI1Z2_SP_L1D3PHI1Z2_L2D3PHI1Z2;
wire TE_L1D3PHI1Z2_L2D3PHI1Z2_SP_L1D3PHI1Z2_L2D3PHI1Z2_wr_en;
wire [5:0] SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1Z2_L2D3PHI1Z2(
.data_in(TE_L1D3PHI1Z2_L2D3PHI1Z2_SP_L1D3PHI1Z2_L2D3PHI1Z2),
.enable(TE_L1D3PHI1Z2_L2D3PHI1Z2_SP_L1D3PHI1Z2_L2D3PHI1Z2_wr_en),
.number_out(SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z2_L2D3PHI2Z2_SP_L1D3PHI1Z2_L2D3PHI2Z2;
wire TE_L1D3PHI1Z2_L2D3PHI2Z2_SP_L1D3PHI1Z2_L2D3PHI2Z2_wr_en;
wire [5:0] SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1Z2_L2D3PHI2Z2(
.data_in(TE_L1D3PHI1Z2_L2D3PHI2Z2_SP_L1D3PHI1Z2_L2D3PHI2Z2),
.enable(TE_L1D3PHI1Z2_L2D3PHI2Z2_SP_L1D3PHI1Z2_L2D3PHI2Z2_wr_en),
.number_out(SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z2_L2D3PHI2Z2_SP_L1D3PHI2Z2_L2D3PHI2Z2;
wire TE_L1D3PHI2Z2_L2D3PHI2Z2_SP_L1D3PHI2Z2_L2D3PHI2Z2_wr_en;
wire [5:0] SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2Z2_L2D3PHI2Z2(
.data_in(TE_L1D3PHI2Z2_L2D3PHI2Z2_SP_L1D3PHI2Z2_L2D3PHI2Z2),
.enable(TE_L1D3PHI2Z2_L2D3PHI2Z2_SP_L1D3PHI2Z2_L2D3PHI2Z2_wr_en),
.number_out(SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z2_L2D3PHI3Z2_SP_L1D3PHI2Z2_L2D3PHI3Z2;
wire TE_L1D3PHI2Z2_L2D3PHI3Z2_SP_L1D3PHI2Z2_L2D3PHI3Z2_wr_en;
wire [5:0] SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2Z2_L2D3PHI3Z2(
.data_in(TE_L1D3PHI2Z2_L2D3PHI3Z2_SP_L1D3PHI2Z2_L2D3PHI3Z2),
.enable(TE_L1D3PHI2Z2_L2D3PHI3Z2_SP_L1D3PHI2Z2_L2D3PHI3Z2_wr_en),
.number_out(SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z2_L2D3PHI3Z2_SP_L1D3PHI3Z2_L2D3PHI3Z2;
wire TE_L1D3PHI3Z2_L2D3PHI3Z2_SP_L1D3PHI3Z2_L2D3PHI3Z2_wr_en;
wire [5:0] SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3Z2_L2D3PHI3Z2(
.data_in(TE_L1D3PHI3Z2_L2D3PHI3Z2_SP_L1D3PHI3Z2_L2D3PHI3Z2),
.enable(TE_L1D3PHI3Z2_L2D3PHI3Z2_SP_L1D3PHI3Z2_L2D3PHI3Z2_wr_en),
.number_out(SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z2_L2D3PHI4Z2_SP_L1D3PHI3Z2_L2D3PHI4Z2;
wire TE_L1D3PHI3Z2_L2D3PHI4Z2_SP_L1D3PHI3Z2_L2D3PHI4Z2_wr_en;
wire [5:0] SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3Z2_L2D3PHI4Z2(
.data_in(TE_L1D3PHI3Z2_L2D3PHI4Z2_SP_L1D3PHI3Z2_L2D3PHI4Z2),
.enable(TE_L1D3PHI3Z2_L2D3PHI4Z2_SP_L1D3PHI3Z2_L2D3PHI4Z2_wr_en),
.number_out(SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L1D3_AS_L1D3n1;
wire VMR_L1D3_AS_L1D3n1_wr_en;
wire [10:0] AS_L1D3n1_TC_L1D3L2D3_read_add;
wire [35:0] AS_L1D3n1_TC_L1D3L2D3;
AllStubs  AS_L1D3n1(
.data_in(VMR_L1D3_AS_L1D3n1),
.enable(VMR_L1D3_AS_L1D3n1_wr_en),
.read_add(AS_L1D3n1_TC_L1D3L2D3_read_add),
.data_out(AS_L1D3n1_TC_L1D3L2D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L2D3_AS_L2D3n1;
wire VMR_L2D3_AS_L2D3n1_wr_en;
wire [10:0] AS_L2D3n1_TC_L1D3L2D3_read_add;
wire [35:0] AS_L2D3n1_TC_L1D3L2D3;
AllStubs  AS_L2D3n1(
.data_in(VMR_L2D3_AS_L2D3n1),
.enable(VMR_L2D3_AS_L2D3n1_wr_en),
.read_add(AS_L2D3n1_TC_L1D3L2D3_read_add),
.data_out(AS_L2D3n1_TC_L1D3L2D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z1_L2D4PHI1Z1_SP_L1D3PHI1Z1_L2D4PHI1Z1;
wire TE_L1D3PHI1Z1_L2D4PHI1Z1_SP_L1D3PHI1Z1_L2D4PHI1Z1_wr_en;
wire [5:0] SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1Z1_L2D4PHI1Z1(
.data_in(TE_L1D3PHI1Z1_L2D4PHI1Z1_SP_L1D3PHI1Z1_L2D4PHI1Z1),
.enable(TE_L1D3PHI1Z1_L2D4PHI1Z1_SP_L1D3PHI1Z1_L2D4PHI1Z1_wr_en),
.number_out(SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z1_L2D4PHI2Z1_SP_L1D3PHI1Z1_L2D4PHI2Z1;
wire TE_L1D3PHI1Z1_L2D4PHI2Z1_SP_L1D3PHI1Z1_L2D4PHI2Z1_wr_en;
wire [5:0] SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1Z1_L2D4PHI2Z1(
.data_in(TE_L1D3PHI1Z1_L2D4PHI2Z1_SP_L1D3PHI1Z1_L2D4PHI2Z1),
.enable(TE_L1D3PHI1Z1_L2D4PHI2Z1_SP_L1D3PHI1Z1_L2D4PHI2Z1_wr_en),
.number_out(SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z1_L2D4PHI2Z1_SP_L1D3PHI2Z1_L2D4PHI2Z1;
wire TE_L1D3PHI2Z1_L2D4PHI2Z1_SP_L1D3PHI2Z1_L2D4PHI2Z1_wr_en;
wire [5:0] SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2Z1_L2D4PHI2Z1(
.data_in(TE_L1D3PHI2Z1_L2D4PHI2Z1_SP_L1D3PHI2Z1_L2D4PHI2Z1),
.enable(TE_L1D3PHI2Z1_L2D4PHI2Z1_SP_L1D3PHI2Z1_L2D4PHI2Z1_wr_en),
.number_out(SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z1_L2D4PHI3Z1_SP_L1D3PHI2Z1_L2D4PHI3Z1;
wire TE_L1D3PHI2Z1_L2D4PHI3Z1_SP_L1D3PHI2Z1_L2D4PHI3Z1_wr_en;
wire [5:0] SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2Z1_L2D4PHI3Z1(
.data_in(TE_L1D3PHI2Z1_L2D4PHI3Z1_SP_L1D3PHI2Z1_L2D4PHI3Z1),
.enable(TE_L1D3PHI2Z1_L2D4PHI3Z1_SP_L1D3PHI2Z1_L2D4PHI3Z1_wr_en),
.number_out(SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z1_L2D4PHI3Z1_SP_L1D3PHI3Z1_L2D4PHI3Z1;
wire TE_L1D3PHI3Z1_L2D4PHI3Z1_SP_L1D3PHI3Z1_L2D4PHI3Z1_wr_en;
wire [5:0] SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3Z1_L2D4PHI3Z1(
.data_in(TE_L1D3PHI3Z1_L2D4PHI3Z1_SP_L1D3PHI3Z1_L2D4PHI3Z1),
.enable(TE_L1D3PHI3Z1_L2D4PHI3Z1_SP_L1D3PHI3Z1_L2D4PHI3Z1_wr_en),
.number_out(SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z1_L2D4PHI4Z1_SP_L1D3PHI3Z1_L2D4PHI4Z1;
wire TE_L1D3PHI3Z1_L2D4PHI4Z1_SP_L1D3PHI3Z1_L2D4PHI4Z1_wr_en;
wire [5:0] SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3Z1_L2D4PHI4Z1(
.data_in(TE_L1D3PHI3Z1_L2D4PHI4Z1_SP_L1D3PHI3Z1_L2D4PHI4Z1),
.enable(TE_L1D3PHI3Z1_L2D4PHI4Z1_SP_L1D3PHI3Z1_L2D4PHI4Z1_wr_en),
.number_out(SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z2_L2D4PHI1Z1_SP_L1D3PHI1Z2_L2D4PHI1Z1;
wire TE_L1D3PHI1Z2_L2D4PHI1Z1_SP_L1D3PHI1Z2_L2D4PHI1Z1_wr_en;
wire [5:0] SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1Z2_L2D4PHI1Z1(
.data_in(TE_L1D3PHI1Z2_L2D4PHI1Z1_SP_L1D3PHI1Z2_L2D4PHI1Z1),
.enable(TE_L1D3PHI1Z2_L2D4PHI1Z1_SP_L1D3PHI1Z2_L2D4PHI1Z1_wr_en),
.number_out(SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z2_L2D4PHI2Z1_SP_L1D3PHI1Z2_L2D4PHI2Z1;
wire TE_L1D3PHI1Z2_L2D4PHI2Z1_SP_L1D3PHI1Z2_L2D4PHI2Z1_wr_en;
wire [5:0] SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1Z2_L2D4PHI2Z1(
.data_in(TE_L1D3PHI1Z2_L2D4PHI2Z1_SP_L1D3PHI1Z2_L2D4PHI2Z1),
.enable(TE_L1D3PHI1Z2_L2D4PHI2Z1_SP_L1D3PHI1Z2_L2D4PHI2Z1_wr_en),
.number_out(SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z2_L2D4PHI2Z1_SP_L1D3PHI2Z2_L2D4PHI2Z1;
wire TE_L1D3PHI2Z2_L2D4PHI2Z1_SP_L1D3PHI2Z2_L2D4PHI2Z1_wr_en;
wire [5:0] SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2Z2_L2D4PHI2Z1(
.data_in(TE_L1D3PHI2Z2_L2D4PHI2Z1_SP_L1D3PHI2Z2_L2D4PHI2Z1),
.enable(TE_L1D3PHI2Z2_L2D4PHI2Z1_SP_L1D3PHI2Z2_L2D4PHI2Z1_wr_en),
.number_out(SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z2_L2D4PHI3Z1_SP_L1D3PHI2Z2_L2D4PHI3Z1;
wire TE_L1D3PHI2Z2_L2D4PHI3Z1_SP_L1D3PHI2Z2_L2D4PHI3Z1_wr_en;
wire [5:0] SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2Z2_L2D4PHI3Z1(
.data_in(TE_L1D3PHI2Z2_L2D4PHI3Z1_SP_L1D3PHI2Z2_L2D4PHI3Z1),
.enable(TE_L1D3PHI2Z2_L2D4PHI3Z1_SP_L1D3PHI2Z2_L2D4PHI3Z1_wr_en),
.number_out(SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z2_L2D4PHI3Z1_SP_L1D3PHI3Z2_L2D4PHI3Z1;
wire TE_L1D3PHI3Z2_L2D4PHI3Z1_SP_L1D3PHI3Z2_L2D4PHI3Z1_wr_en;
wire [5:0] SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3Z2_L2D4PHI3Z1(
.data_in(TE_L1D3PHI3Z2_L2D4PHI3Z1_SP_L1D3PHI3Z2_L2D4PHI3Z1),
.enable(TE_L1D3PHI3Z2_L2D4PHI3Z1_SP_L1D3PHI3Z2_L2D4PHI3Z1_wr_en),
.number_out(SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z2_L2D4PHI4Z1_SP_L1D3PHI3Z2_L2D4PHI4Z1;
wire TE_L1D3PHI3Z2_L2D4PHI4Z1_SP_L1D3PHI3Z2_L2D4PHI4Z1_wr_en;
wire [5:0] SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3Z2_L2D4PHI4Z1(
.data_in(TE_L1D3PHI3Z2_L2D4PHI4Z1_SP_L1D3PHI3Z2_L2D4PHI4Z1),
.enable(TE_L1D3PHI3Z2_L2D4PHI4Z1_SP_L1D3PHI3Z2_L2D4PHI4Z1_wr_en),
.number_out(SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z2_L2D4PHI1Z2_SP_L1D3PHI1Z2_L2D4PHI1Z2;
wire TE_L1D3PHI1Z2_L2D4PHI1Z2_SP_L1D3PHI1Z2_L2D4PHI1Z2_wr_en;
wire [5:0] SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1Z2_L2D4PHI1Z2(
.data_in(TE_L1D3PHI1Z2_L2D4PHI1Z2_SP_L1D3PHI1Z2_L2D4PHI1Z2),
.enable(TE_L1D3PHI1Z2_L2D4PHI1Z2_SP_L1D3PHI1Z2_L2D4PHI1Z2_wr_en),
.number_out(SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI1Z2_L2D4PHI2Z2_SP_L1D3PHI1Z2_L2D4PHI2Z2;
wire TE_L1D3PHI1Z2_L2D4PHI2Z2_SP_L1D3PHI1Z2_L2D4PHI2Z2_wr_en;
wire [5:0] SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1Z2_L2D4PHI2Z2(
.data_in(TE_L1D3PHI1Z2_L2D4PHI2Z2_SP_L1D3PHI1Z2_L2D4PHI2Z2),
.enable(TE_L1D3PHI1Z2_L2D4PHI2Z2_SP_L1D3PHI1Z2_L2D4PHI2Z2_wr_en),
.number_out(SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z2_L2D4PHI2Z2_SP_L1D3PHI2Z2_L2D4PHI2Z2;
wire TE_L1D3PHI2Z2_L2D4PHI2Z2_SP_L1D3PHI2Z2_L2D4PHI2Z2_wr_en;
wire [5:0] SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2Z2_L2D4PHI2Z2(
.data_in(TE_L1D3PHI2Z2_L2D4PHI2Z2_SP_L1D3PHI2Z2_L2D4PHI2Z2),
.enable(TE_L1D3PHI2Z2_L2D4PHI2Z2_SP_L1D3PHI2Z2_L2D4PHI2Z2_wr_en),
.number_out(SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI2Z2_L2D4PHI3Z2_SP_L1D3PHI2Z2_L2D4PHI3Z2;
wire TE_L1D3PHI2Z2_L2D4PHI3Z2_SP_L1D3PHI2Z2_L2D4PHI3Z2_wr_en;
wire [5:0] SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2Z2_L2D4PHI3Z2(
.data_in(TE_L1D3PHI2Z2_L2D4PHI3Z2_SP_L1D3PHI2Z2_L2D4PHI3Z2),
.enable(TE_L1D3PHI2Z2_L2D4PHI3Z2_SP_L1D3PHI2Z2_L2D4PHI3Z2_wr_en),
.number_out(SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z2_L2D4PHI3Z2_SP_L1D3PHI3Z2_L2D4PHI3Z2;
wire TE_L1D3PHI3Z2_L2D4PHI3Z2_SP_L1D3PHI3Z2_L2D4PHI3Z2_wr_en;
wire [5:0] SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3Z2_L2D4PHI3Z2(
.data_in(TE_L1D3PHI3Z2_L2D4PHI3Z2_SP_L1D3PHI3Z2_L2D4PHI3Z2),
.enable(TE_L1D3PHI3Z2_L2D4PHI3Z2_SP_L1D3PHI3Z2_L2D4PHI3Z2_wr_en),
.number_out(SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D3PHI3Z2_L2D4PHI4Z2_SP_L1D3PHI3Z2_L2D4PHI4Z2;
wire TE_L1D3PHI3Z2_L2D4PHI4Z2_SP_L1D3PHI3Z2_L2D4PHI4Z2_wr_en;
wire [5:0] SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3Z2_L2D4PHI4Z2(
.data_in(TE_L1D3PHI3Z2_L2D4PHI4Z2_SP_L1D3PHI3Z2_L2D4PHI4Z2),
.enable(TE_L1D3PHI3Z2_L2D4PHI4Z2_SP_L1D3PHI3Z2_L2D4PHI4Z2_wr_en),
.number_out(SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L1D3_AS_L1D3n2;
wire VMR_L1D3_AS_L1D3n2_wr_en;
wire [10:0] AS_L1D3n2_TC_L1D3L2D4_read_add;
wire [35:0] AS_L1D3n2_TC_L1D3L2D4;
AllStubs  AS_L1D3n2(
.data_in(VMR_L1D3_AS_L1D3n2),
.enable(VMR_L1D3_AS_L1D3n2_wr_en),
.read_add(AS_L1D3n2_TC_L1D3L2D4_read_add),
.data_out(AS_L1D3n2_TC_L1D3L2D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L2D4_AS_L2D4n1;
wire VMR_L2D4_AS_L2D4n1_wr_en;
wire [10:0] AS_L2D4n1_TC_L1D3L2D4_read_add;
wire [35:0] AS_L2D4n1_TC_L1D3L2D4;
AllStubs  AS_L2D4n1(
.data_in(VMR_L2D4_AS_L2D4n1),
.enable(VMR_L2D4_AS_L2D4n1_wr_en),
.read_add(AS_L2D4n1_TC_L1D3L2D4_read_add),
.data_out(AS_L2D4n1_TC_L1D3L2D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D4PHI1Z1_L2D4PHI1Z2_SP_L1D4PHI1Z1_L2D4PHI1Z2;
wire TE_L1D4PHI1Z1_L2D4PHI1Z2_SP_L1D4PHI1Z1_L2D4PHI1Z2_wr_en;
wire [5:0] SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI1Z1_L2D4PHI1Z2(
.data_in(TE_L1D4PHI1Z1_L2D4PHI1Z2_SP_L1D4PHI1Z1_L2D4PHI1Z2),
.enable(TE_L1D4PHI1Z1_L2D4PHI1Z2_SP_L1D4PHI1Z1_L2D4PHI1Z2_wr_en),
.number_out(SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D4PHI1Z1_L2D4PHI2Z2_SP_L1D4PHI1Z1_L2D4PHI2Z2;
wire TE_L1D4PHI1Z1_L2D4PHI2Z2_SP_L1D4PHI1Z1_L2D4PHI2Z2_wr_en;
wire [5:0] SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI1Z1_L2D4PHI2Z2(
.data_in(TE_L1D4PHI1Z1_L2D4PHI2Z2_SP_L1D4PHI1Z1_L2D4PHI2Z2),
.enable(TE_L1D4PHI1Z1_L2D4PHI2Z2_SP_L1D4PHI1Z1_L2D4PHI2Z2_wr_en),
.number_out(SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D4PHI2Z1_L2D4PHI2Z2_SP_L1D4PHI2Z1_L2D4PHI2Z2;
wire TE_L1D4PHI2Z1_L2D4PHI2Z2_SP_L1D4PHI2Z1_L2D4PHI2Z2_wr_en;
wire [5:0] SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI2Z1_L2D4PHI2Z2(
.data_in(TE_L1D4PHI2Z1_L2D4PHI2Z2_SP_L1D4PHI2Z1_L2D4PHI2Z2),
.enable(TE_L1D4PHI2Z1_L2D4PHI2Z2_SP_L1D4PHI2Z1_L2D4PHI2Z2_wr_en),
.number_out(SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D4PHI2Z1_L2D4PHI3Z2_SP_L1D4PHI2Z1_L2D4PHI3Z2;
wire TE_L1D4PHI2Z1_L2D4PHI3Z2_SP_L1D4PHI2Z1_L2D4PHI3Z2_wr_en;
wire [5:0] SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI2Z1_L2D4PHI3Z2(
.data_in(TE_L1D4PHI2Z1_L2D4PHI3Z2_SP_L1D4PHI2Z1_L2D4PHI3Z2),
.enable(TE_L1D4PHI2Z1_L2D4PHI3Z2_SP_L1D4PHI2Z1_L2D4PHI3Z2_wr_en),
.number_out(SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D4PHI3Z1_L2D4PHI3Z2_SP_L1D4PHI3Z1_L2D4PHI3Z2;
wire TE_L1D4PHI3Z1_L2D4PHI3Z2_SP_L1D4PHI3Z1_L2D4PHI3Z2_wr_en;
wire [5:0] SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI3Z1_L2D4PHI3Z2(
.data_in(TE_L1D4PHI3Z1_L2D4PHI3Z2_SP_L1D4PHI3Z1_L2D4PHI3Z2),
.enable(TE_L1D4PHI3Z1_L2D4PHI3Z2_SP_L1D4PHI3Z1_L2D4PHI3Z2_wr_en),
.number_out(SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L1D4PHI3Z1_L2D4PHI4Z2_SP_L1D4PHI3Z1_L2D4PHI4Z2;
wire TE_L1D4PHI3Z1_L2D4PHI4Z2_SP_L1D4PHI3Z1_L2D4PHI4Z2_wr_en;
wire [5:0] SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI3Z1_L2D4PHI4Z2(
.data_in(TE_L1D4PHI3Z1_L2D4PHI4Z2_SP_L1D4PHI3Z1_L2D4PHI4Z2),
.enable(TE_L1D4PHI3Z1_L2D4PHI4Z2_SP_L1D4PHI3Z1_L2D4PHI4Z2_wr_en),
.number_out(SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L1D4_AS_L1D4n1;
wire VMR_L1D4_AS_L1D4n1_wr_en;
wire [10:0] AS_L1D4n1_TC_L1D4L2D4_read_add;
wire [35:0] AS_L1D4n1_TC_L1D4L2D4;
AllStubs  AS_L1D4n1(
.data_in(VMR_L1D4_AS_L1D4n1),
.enable(VMR_L1D4_AS_L1D4n1_wr_en),
.read_add(AS_L1D4n1_TC_L1D4L2D4_read_add),
.data_out(AS_L1D4n1_TC_L1D4L2D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L2D4_AS_L2D4n2;
wire VMR_L2D4_AS_L2D4n2_wr_en;
wire [10:0] AS_L2D4n2_TC_L1D4L2D4_read_add;
wire [35:0] AS_L2D4n2_TC_L1D4L2D4;
AllStubs  AS_L2D4n2(
.data_in(VMR_L2D4_AS_L2D4n2),
.enable(VMR_L2D4_AS_L2D4n2_wr_en),
.read_add(AS_L2D4n2_TC_L1D4L2D4_read_add),
.data_out(AS_L2D4n2_TC_L1D4L2D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI1Z1_L4D3PHI1Z1_SP_L3D3PHI1Z1_L4D3PHI1Z1;
wire TE_L3D3PHI1Z1_L4D3PHI1Z1_SP_L3D3PHI1Z1_L4D3PHI1Z1_wr_en;
wire [5:0] SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1Z1_L4D3PHI1Z1(
.data_in(TE_L3D3PHI1Z1_L4D3PHI1Z1_SP_L3D3PHI1Z1_L4D3PHI1Z1),
.enable(TE_L3D3PHI1Z1_L4D3PHI1Z1_SP_L3D3PHI1Z1_L4D3PHI1Z1_wr_en),
.number_out(SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI1Z1_L4D3PHI2Z1_SP_L3D3PHI1Z1_L4D3PHI2Z1;
wire TE_L3D3PHI1Z1_L4D3PHI2Z1_SP_L3D3PHI1Z1_L4D3PHI2Z1_wr_en;
wire [5:0] SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1Z1_L4D3PHI2Z1(
.data_in(TE_L3D3PHI1Z1_L4D3PHI2Z1_SP_L3D3PHI1Z1_L4D3PHI2Z1),
.enable(TE_L3D3PHI1Z1_L4D3PHI2Z1_SP_L3D3PHI1Z1_L4D3PHI2Z1_wr_en),
.number_out(SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI2Z1_L4D3PHI2Z1_SP_L3D3PHI2Z1_L4D3PHI2Z1;
wire TE_L3D3PHI2Z1_L4D3PHI2Z1_SP_L3D3PHI2Z1_L4D3PHI2Z1_wr_en;
wire [5:0] SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2Z1_L4D3PHI2Z1(
.data_in(TE_L3D3PHI2Z1_L4D3PHI2Z1_SP_L3D3PHI2Z1_L4D3PHI2Z1),
.enable(TE_L3D3PHI2Z1_L4D3PHI2Z1_SP_L3D3PHI2Z1_L4D3PHI2Z1_wr_en),
.number_out(SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI2Z1_L4D3PHI3Z1_SP_L3D3PHI2Z1_L4D3PHI3Z1;
wire TE_L3D3PHI2Z1_L4D3PHI3Z1_SP_L3D3PHI2Z1_L4D3PHI3Z1_wr_en;
wire [5:0] SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2Z1_L4D3PHI3Z1(
.data_in(TE_L3D3PHI2Z1_L4D3PHI3Z1_SP_L3D3PHI2Z1_L4D3PHI3Z1),
.enable(TE_L3D3PHI2Z1_L4D3PHI3Z1_SP_L3D3PHI2Z1_L4D3PHI3Z1_wr_en),
.number_out(SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI3Z1_L4D3PHI3Z1_SP_L3D3PHI3Z1_L4D3PHI3Z1;
wire TE_L3D3PHI3Z1_L4D3PHI3Z1_SP_L3D3PHI3Z1_L4D3PHI3Z1_wr_en;
wire [5:0] SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3Z1_L4D3PHI3Z1(
.data_in(TE_L3D3PHI3Z1_L4D3PHI3Z1_SP_L3D3PHI3Z1_L4D3PHI3Z1),
.enable(TE_L3D3PHI3Z1_L4D3PHI3Z1_SP_L3D3PHI3Z1_L4D3PHI3Z1_wr_en),
.number_out(SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI3Z1_L4D3PHI4Z1_SP_L3D3PHI3Z1_L4D3PHI4Z1;
wire TE_L3D3PHI3Z1_L4D3PHI4Z1_SP_L3D3PHI3Z1_L4D3PHI4Z1_wr_en;
wire [5:0] SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3Z1_L4D3PHI4Z1(
.data_in(TE_L3D3PHI3Z1_L4D3PHI4Z1_SP_L3D3PHI3Z1_L4D3PHI4Z1),
.enable(TE_L3D3PHI3Z1_L4D3PHI4Z1_SP_L3D3PHI3Z1_L4D3PHI4Z1_wr_en),
.number_out(SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI1Z1_L4D3PHI1Z2_SP_L3D3PHI1Z1_L4D3PHI1Z2;
wire TE_L3D3PHI1Z1_L4D3PHI1Z2_SP_L3D3PHI1Z1_L4D3PHI1Z2_wr_en;
wire [5:0] SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1Z1_L4D3PHI1Z2(
.data_in(TE_L3D3PHI1Z1_L4D3PHI1Z2_SP_L3D3PHI1Z1_L4D3PHI1Z2),
.enable(TE_L3D3PHI1Z1_L4D3PHI1Z2_SP_L3D3PHI1Z1_L4D3PHI1Z2_wr_en),
.number_out(SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI1Z1_L4D3PHI2Z2_SP_L3D3PHI1Z1_L4D3PHI2Z2;
wire TE_L3D3PHI1Z1_L4D3PHI2Z2_SP_L3D3PHI1Z1_L4D3PHI2Z2_wr_en;
wire [5:0] SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1Z1_L4D3PHI2Z2(
.data_in(TE_L3D3PHI1Z1_L4D3PHI2Z2_SP_L3D3PHI1Z1_L4D3PHI2Z2),
.enable(TE_L3D3PHI1Z1_L4D3PHI2Z2_SP_L3D3PHI1Z1_L4D3PHI2Z2_wr_en),
.number_out(SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI2Z1_L4D3PHI2Z2_SP_L3D3PHI2Z1_L4D3PHI2Z2;
wire TE_L3D3PHI2Z1_L4D3PHI2Z2_SP_L3D3PHI2Z1_L4D3PHI2Z2_wr_en;
wire [5:0] SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2Z1_L4D3PHI2Z2(
.data_in(TE_L3D3PHI2Z1_L4D3PHI2Z2_SP_L3D3PHI2Z1_L4D3PHI2Z2),
.enable(TE_L3D3PHI2Z1_L4D3PHI2Z2_SP_L3D3PHI2Z1_L4D3PHI2Z2_wr_en),
.number_out(SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI2Z1_L4D3PHI3Z2_SP_L3D3PHI2Z1_L4D3PHI3Z2;
wire TE_L3D3PHI2Z1_L4D3PHI3Z2_SP_L3D3PHI2Z1_L4D3PHI3Z2_wr_en;
wire [5:0] SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2Z1_L4D3PHI3Z2(
.data_in(TE_L3D3PHI2Z1_L4D3PHI3Z2_SP_L3D3PHI2Z1_L4D3PHI3Z2),
.enable(TE_L3D3PHI2Z1_L4D3PHI3Z2_SP_L3D3PHI2Z1_L4D3PHI3Z2_wr_en),
.number_out(SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI3Z1_L4D3PHI3Z2_SP_L3D3PHI3Z1_L4D3PHI3Z2;
wire TE_L3D3PHI3Z1_L4D3PHI3Z2_SP_L3D3PHI3Z1_L4D3PHI3Z2_wr_en;
wire [5:0] SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3Z1_L4D3PHI3Z2(
.data_in(TE_L3D3PHI3Z1_L4D3PHI3Z2_SP_L3D3PHI3Z1_L4D3PHI3Z2),
.enable(TE_L3D3PHI3Z1_L4D3PHI3Z2_SP_L3D3PHI3Z1_L4D3PHI3Z2_wr_en),
.number_out(SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI3Z1_L4D3PHI4Z2_SP_L3D3PHI3Z1_L4D3PHI4Z2;
wire TE_L3D3PHI3Z1_L4D3PHI4Z2_SP_L3D3PHI3Z1_L4D3PHI4Z2_wr_en;
wire [5:0] SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3Z1_L4D3PHI4Z2(
.data_in(TE_L3D3PHI3Z1_L4D3PHI4Z2_SP_L3D3PHI3Z1_L4D3PHI4Z2),
.enable(TE_L3D3PHI3Z1_L4D3PHI4Z2_SP_L3D3PHI3Z1_L4D3PHI4Z2_wr_en),
.number_out(SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI1Z2_L4D3PHI1Z2_SP_L3D3PHI1Z2_L4D3PHI1Z2;
wire TE_L3D3PHI1Z2_L4D3PHI1Z2_SP_L3D3PHI1Z2_L4D3PHI1Z2_wr_en;
wire [5:0] SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1Z2_L4D3PHI1Z2(
.data_in(TE_L3D3PHI1Z2_L4D3PHI1Z2_SP_L3D3PHI1Z2_L4D3PHI1Z2),
.enable(TE_L3D3PHI1Z2_L4D3PHI1Z2_SP_L3D3PHI1Z2_L4D3PHI1Z2_wr_en),
.number_out(SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI1Z2_L4D3PHI2Z2_SP_L3D3PHI1Z2_L4D3PHI2Z2;
wire TE_L3D3PHI1Z2_L4D3PHI2Z2_SP_L3D3PHI1Z2_L4D3PHI2Z2_wr_en;
wire [5:0] SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1Z2_L4D3PHI2Z2(
.data_in(TE_L3D3PHI1Z2_L4D3PHI2Z2_SP_L3D3PHI1Z2_L4D3PHI2Z2),
.enable(TE_L3D3PHI1Z2_L4D3PHI2Z2_SP_L3D3PHI1Z2_L4D3PHI2Z2_wr_en),
.number_out(SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI2Z2_L4D3PHI2Z2_SP_L3D3PHI2Z2_L4D3PHI2Z2;
wire TE_L3D3PHI2Z2_L4D3PHI2Z2_SP_L3D3PHI2Z2_L4D3PHI2Z2_wr_en;
wire [5:0] SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2Z2_L4D3PHI2Z2(
.data_in(TE_L3D3PHI2Z2_L4D3PHI2Z2_SP_L3D3PHI2Z2_L4D3PHI2Z2),
.enable(TE_L3D3PHI2Z2_L4D3PHI2Z2_SP_L3D3PHI2Z2_L4D3PHI2Z2_wr_en),
.number_out(SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI2Z2_L4D3PHI3Z2_SP_L3D3PHI2Z2_L4D3PHI3Z2;
wire TE_L3D3PHI2Z2_L4D3PHI3Z2_SP_L3D3PHI2Z2_L4D3PHI3Z2_wr_en;
wire [5:0] SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2Z2_L4D3PHI3Z2(
.data_in(TE_L3D3PHI2Z2_L4D3PHI3Z2_SP_L3D3PHI2Z2_L4D3PHI3Z2),
.enable(TE_L3D3PHI2Z2_L4D3PHI3Z2_SP_L3D3PHI2Z2_L4D3PHI3Z2_wr_en),
.number_out(SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI3Z2_L4D3PHI3Z2_SP_L3D3PHI3Z2_L4D3PHI3Z2;
wire TE_L3D3PHI3Z2_L4D3PHI3Z2_SP_L3D3PHI3Z2_L4D3PHI3Z2_wr_en;
wire [5:0] SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3Z2_L4D3PHI3Z2(
.data_in(TE_L3D3PHI3Z2_L4D3PHI3Z2_SP_L3D3PHI3Z2_L4D3PHI3Z2),
.enable(TE_L3D3PHI3Z2_L4D3PHI3Z2_SP_L3D3PHI3Z2_L4D3PHI3Z2_wr_en),
.number_out(SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI3Z2_L4D3PHI4Z2_SP_L3D3PHI3Z2_L4D3PHI4Z2;
wire TE_L3D3PHI3Z2_L4D3PHI4Z2_SP_L3D3PHI3Z2_L4D3PHI4Z2_wr_en;
wire [5:0] SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3Z2_L4D3PHI4Z2(
.data_in(TE_L3D3PHI3Z2_L4D3PHI4Z2_SP_L3D3PHI3Z2_L4D3PHI4Z2),
.enable(TE_L3D3PHI3Z2_L4D3PHI4Z2_SP_L3D3PHI3Z2_L4D3PHI4Z2_wr_en),
.number_out(SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L3D3_AS_L3D3n1;
wire VMR_L3D3_AS_L3D3n1_wr_en;
wire [10:0] AS_L3D3n1_TC_L3D3L4D3_read_add;
wire [35:0] AS_L3D3n1_TC_L3D3L4D3;
AllStubs  AS_L3D3n1(
.data_in(VMR_L3D3_AS_L3D3n1),
.enable(VMR_L3D3_AS_L3D3n1_wr_en),
.read_add(AS_L3D3n1_TC_L3D3L4D3_read_add),
.data_out(AS_L3D3n1_TC_L3D3L4D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L4D3_AS_L4D3n1;
wire VMR_L4D3_AS_L4D3n1_wr_en;
wire [10:0] AS_L4D3n1_TC_L3D3L4D3_read_add;
wire [35:0] AS_L4D3n1_TC_L3D3L4D3;
AllStubs  AS_L4D3n1(
.data_in(VMR_L4D3_AS_L4D3n1),
.enable(VMR_L4D3_AS_L4D3n1_wr_en),
.read_add(AS_L4D3n1_TC_L3D3L4D3_read_add),
.data_out(AS_L4D3n1_TC_L3D3L4D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI1Z2_L4D4PHI1Z1_SP_L3D3PHI1Z2_L4D4PHI1Z1;
wire TE_L3D3PHI1Z2_L4D4PHI1Z1_SP_L3D3PHI1Z2_L4D4PHI1Z1_wr_en;
wire [5:0] SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI1Z2_L4D4PHI1Z1(
.data_in(TE_L3D3PHI1Z2_L4D4PHI1Z1_SP_L3D3PHI1Z2_L4D4PHI1Z1),
.enable(TE_L3D3PHI1Z2_L4D4PHI1Z1_SP_L3D3PHI1Z2_L4D4PHI1Z1_wr_en),
.number_out(SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI1Z2_L4D4PHI2Z1_SP_L3D3PHI1Z2_L4D4PHI2Z1;
wire TE_L3D3PHI1Z2_L4D4PHI2Z1_SP_L3D3PHI1Z2_L4D4PHI2Z1_wr_en;
wire [5:0] SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI1Z2_L4D4PHI2Z1(
.data_in(TE_L3D3PHI1Z2_L4D4PHI2Z1_SP_L3D3PHI1Z2_L4D4PHI2Z1),
.enable(TE_L3D3PHI1Z2_L4D4PHI2Z1_SP_L3D3PHI1Z2_L4D4PHI2Z1_wr_en),
.number_out(SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI2Z2_L4D4PHI2Z1_SP_L3D3PHI2Z2_L4D4PHI2Z1;
wire TE_L3D3PHI2Z2_L4D4PHI2Z1_SP_L3D3PHI2Z2_L4D4PHI2Z1_wr_en;
wire [5:0] SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI2Z2_L4D4PHI2Z1(
.data_in(TE_L3D3PHI2Z2_L4D4PHI2Z1_SP_L3D3PHI2Z2_L4D4PHI2Z1),
.enable(TE_L3D3PHI2Z2_L4D4PHI2Z1_SP_L3D3PHI2Z2_L4D4PHI2Z1_wr_en),
.number_out(SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI2Z2_L4D4PHI3Z1_SP_L3D3PHI2Z2_L4D4PHI3Z1;
wire TE_L3D3PHI2Z2_L4D4PHI3Z1_SP_L3D3PHI2Z2_L4D4PHI3Z1_wr_en;
wire [5:0] SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI2Z2_L4D4PHI3Z1(
.data_in(TE_L3D3PHI2Z2_L4D4PHI3Z1_SP_L3D3PHI2Z2_L4D4PHI3Z1),
.enable(TE_L3D3PHI2Z2_L4D4PHI3Z1_SP_L3D3PHI2Z2_L4D4PHI3Z1_wr_en),
.number_out(SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI3Z2_L4D4PHI3Z1_SP_L3D3PHI3Z2_L4D4PHI3Z1;
wire TE_L3D3PHI3Z2_L4D4PHI3Z1_SP_L3D3PHI3Z2_L4D4PHI3Z1_wr_en;
wire [5:0] SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI3Z2_L4D4PHI3Z1(
.data_in(TE_L3D3PHI3Z2_L4D4PHI3Z1_SP_L3D3PHI3Z2_L4D4PHI3Z1),
.enable(TE_L3D3PHI3Z2_L4D4PHI3Z1_SP_L3D3PHI3Z2_L4D4PHI3Z1_wr_en),
.number_out(SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D3PHI3Z2_L4D4PHI4Z1_SP_L3D3PHI3Z2_L4D4PHI4Z1;
wire TE_L3D3PHI3Z2_L4D4PHI4Z1_SP_L3D3PHI3Z2_L4D4PHI4Z1_wr_en;
wire [5:0] SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI3Z2_L4D4PHI4Z1(
.data_in(TE_L3D3PHI3Z2_L4D4PHI4Z1_SP_L3D3PHI3Z2_L4D4PHI4Z1),
.enable(TE_L3D3PHI3Z2_L4D4PHI4Z1_SP_L3D3PHI3Z2_L4D4PHI4Z1_wr_en),
.number_out(SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L3D3_AS_L3D3n2;
wire VMR_L3D3_AS_L3D3n2_wr_en;
wire [10:0] AS_L3D3n2_TC_L3D3L4D4_read_add;
wire [35:0] AS_L3D3n2_TC_L3D3L4D4;
AllStubs  AS_L3D3n2(
.data_in(VMR_L3D3_AS_L3D3n2),
.enable(VMR_L3D3_AS_L3D3n2_wr_en),
.read_add(AS_L3D3n2_TC_L3D3L4D4_read_add),
.data_out(AS_L3D3n2_TC_L3D3L4D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L4D4_AS_L4D4n1;
wire VMR_L4D4_AS_L4D4n1_wr_en;
wire [10:0] AS_L4D4n1_TC_L3D3L4D4_read_add;
wire [35:0] AS_L4D4n1_TC_L3D3L4D4;
AllStubs  AS_L4D4n1(
.data_in(VMR_L4D4_AS_L4D4n1),
.enable(VMR_L4D4_AS_L4D4n1_wr_en),
.read_add(AS_L4D4n1_TC_L3D3L4D4_read_add),
.data_out(AS_L4D4n1_TC_L3D3L4D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI1Z1_L4D4PHI1Z1_SP_L3D4PHI1Z1_L4D4PHI1Z1;
wire TE_L3D4PHI1Z1_L4D4PHI1Z1_SP_L3D4PHI1Z1_L4D4PHI1Z1_wr_en;
wire [5:0] SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1Z1_L4D4PHI1Z1(
.data_in(TE_L3D4PHI1Z1_L4D4PHI1Z1_SP_L3D4PHI1Z1_L4D4PHI1Z1),
.enable(TE_L3D4PHI1Z1_L4D4PHI1Z1_SP_L3D4PHI1Z1_L4D4PHI1Z1_wr_en),
.number_out(SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI1Z1_L4D4PHI2Z1_SP_L3D4PHI1Z1_L4D4PHI2Z1;
wire TE_L3D4PHI1Z1_L4D4PHI2Z1_SP_L3D4PHI1Z1_L4D4PHI2Z1_wr_en;
wire [5:0] SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1Z1_L4D4PHI2Z1(
.data_in(TE_L3D4PHI1Z1_L4D4PHI2Z1_SP_L3D4PHI1Z1_L4D4PHI2Z1),
.enable(TE_L3D4PHI1Z1_L4D4PHI2Z1_SP_L3D4PHI1Z1_L4D4PHI2Z1_wr_en),
.number_out(SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI2Z1_L4D4PHI2Z1_SP_L3D4PHI2Z1_L4D4PHI2Z1;
wire TE_L3D4PHI2Z1_L4D4PHI2Z1_SP_L3D4PHI2Z1_L4D4PHI2Z1_wr_en;
wire [5:0] SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2Z1_L4D4PHI2Z1(
.data_in(TE_L3D4PHI2Z1_L4D4PHI2Z1_SP_L3D4PHI2Z1_L4D4PHI2Z1),
.enable(TE_L3D4PHI2Z1_L4D4PHI2Z1_SP_L3D4PHI2Z1_L4D4PHI2Z1_wr_en),
.number_out(SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI2Z1_L4D4PHI3Z1_SP_L3D4PHI2Z1_L4D4PHI3Z1;
wire TE_L3D4PHI2Z1_L4D4PHI3Z1_SP_L3D4PHI2Z1_L4D4PHI3Z1_wr_en;
wire [5:0] SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2Z1_L4D4PHI3Z1(
.data_in(TE_L3D4PHI2Z1_L4D4PHI3Z1_SP_L3D4PHI2Z1_L4D4PHI3Z1),
.enable(TE_L3D4PHI2Z1_L4D4PHI3Z1_SP_L3D4PHI2Z1_L4D4PHI3Z1_wr_en),
.number_out(SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI3Z1_L4D4PHI3Z1_SP_L3D4PHI3Z1_L4D4PHI3Z1;
wire TE_L3D4PHI3Z1_L4D4PHI3Z1_SP_L3D4PHI3Z1_L4D4PHI3Z1_wr_en;
wire [5:0] SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3Z1_L4D4PHI3Z1(
.data_in(TE_L3D4PHI3Z1_L4D4PHI3Z1_SP_L3D4PHI3Z1_L4D4PHI3Z1),
.enable(TE_L3D4PHI3Z1_L4D4PHI3Z1_SP_L3D4PHI3Z1_L4D4PHI3Z1_wr_en),
.number_out(SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI3Z1_L4D4PHI4Z1_SP_L3D4PHI3Z1_L4D4PHI4Z1;
wire TE_L3D4PHI3Z1_L4D4PHI4Z1_SP_L3D4PHI3Z1_L4D4PHI4Z1_wr_en;
wire [5:0] SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3Z1_L4D4PHI4Z1(
.data_in(TE_L3D4PHI3Z1_L4D4PHI4Z1_SP_L3D4PHI3Z1_L4D4PHI4Z1),
.enable(TE_L3D4PHI3Z1_L4D4PHI4Z1_SP_L3D4PHI3Z1_L4D4PHI4Z1_wr_en),
.number_out(SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI1Z1_L4D4PHI1Z2_SP_L3D4PHI1Z1_L4D4PHI1Z2;
wire TE_L3D4PHI1Z1_L4D4PHI1Z2_SP_L3D4PHI1Z1_L4D4PHI1Z2_wr_en;
wire [5:0] SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1Z1_L4D4PHI1Z2(
.data_in(TE_L3D4PHI1Z1_L4D4PHI1Z2_SP_L3D4PHI1Z1_L4D4PHI1Z2),
.enable(TE_L3D4PHI1Z1_L4D4PHI1Z2_SP_L3D4PHI1Z1_L4D4PHI1Z2_wr_en),
.number_out(SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI1Z1_L4D4PHI2Z2_SP_L3D4PHI1Z1_L4D4PHI2Z2;
wire TE_L3D4PHI1Z1_L4D4PHI2Z2_SP_L3D4PHI1Z1_L4D4PHI2Z2_wr_en;
wire [5:0] SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1Z1_L4D4PHI2Z2(
.data_in(TE_L3D4PHI1Z1_L4D4PHI2Z2_SP_L3D4PHI1Z1_L4D4PHI2Z2),
.enable(TE_L3D4PHI1Z1_L4D4PHI2Z2_SP_L3D4PHI1Z1_L4D4PHI2Z2_wr_en),
.number_out(SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI2Z1_L4D4PHI2Z2_SP_L3D4PHI2Z1_L4D4PHI2Z2;
wire TE_L3D4PHI2Z1_L4D4PHI2Z2_SP_L3D4PHI2Z1_L4D4PHI2Z2_wr_en;
wire [5:0] SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2Z1_L4D4PHI2Z2(
.data_in(TE_L3D4PHI2Z1_L4D4PHI2Z2_SP_L3D4PHI2Z1_L4D4PHI2Z2),
.enable(TE_L3D4PHI2Z1_L4D4PHI2Z2_SP_L3D4PHI2Z1_L4D4PHI2Z2_wr_en),
.number_out(SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI2Z1_L4D4PHI3Z2_SP_L3D4PHI2Z1_L4D4PHI3Z2;
wire TE_L3D4PHI2Z1_L4D4PHI3Z2_SP_L3D4PHI2Z1_L4D4PHI3Z2_wr_en;
wire [5:0] SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2Z1_L4D4PHI3Z2(
.data_in(TE_L3D4PHI2Z1_L4D4PHI3Z2_SP_L3D4PHI2Z1_L4D4PHI3Z2),
.enable(TE_L3D4PHI2Z1_L4D4PHI3Z2_SP_L3D4PHI2Z1_L4D4PHI3Z2_wr_en),
.number_out(SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI3Z1_L4D4PHI3Z2_SP_L3D4PHI3Z1_L4D4PHI3Z2;
wire TE_L3D4PHI3Z1_L4D4PHI3Z2_SP_L3D4PHI3Z1_L4D4PHI3Z2_wr_en;
wire [5:0] SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3Z1_L4D4PHI3Z2(
.data_in(TE_L3D4PHI3Z1_L4D4PHI3Z2_SP_L3D4PHI3Z1_L4D4PHI3Z2),
.enable(TE_L3D4PHI3Z1_L4D4PHI3Z2_SP_L3D4PHI3Z1_L4D4PHI3Z2_wr_en),
.number_out(SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI3Z1_L4D4PHI4Z2_SP_L3D4PHI3Z1_L4D4PHI4Z2;
wire TE_L3D4PHI3Z1_L4D4PHI4Z2_SP_L3D4PHI3Z1_L4D4PHI4Z2_wr_en;
wire [5:0] SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3Z1_L4D4PHI4Z2(
.data_in(TE_L3D4PHI3Z1_L4D4PHI4Z2_SP_L3D4PHI3Z1_L4D4PHI4Z2),
.enable(TE_L3D4PHI3Z1_L4D4PHI4Z2_SP_L3D4PHI3Z1_L4D4PHI4Z2_wr_en),
.number_out(SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI1Z2_L4D4PHI1Z2_SP_L3D4PHI1Z2_L4D4PHI1Z2;
wire TE_L3D4PHI1Z2_L4D4PHI1Z2_SP_L3D4PHI1Z2_L4D4PHI1Z2_wr_en;
wire [5:0] SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1Z2_L4D4PHI1Z2(
.data_in(TE_L3D4PHI1Z2_L4D4PHI1Z2_SP_L3D4PHI1Z2_L4D4PHI1Z2),
.enable(TE_L3D4PHI1Z2_L4D4PHI1Z2_SP_L3D4PHI1Z2_L4D4PHI1Z2_wr_en),
.number_out(SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI1Z2_L4D4PHI2Z2_SP_L3D4PHI1Z2_L4D4PHI2Z2;
wire TE_L3D4PHI1Z2_L4D4PHI2Z2_SP_L3D4PHI1Z2_L4D4PHI2Z2_wr_en;
wire [5:0] SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1Z2_L4D4PHI2Z2(
.data_in(TE_L3D4PHI1Z2_L4D4PHI2Z2_SP_L3D4PHI1Z2_L4D4PHI2Z2),
.enable(TE_L3D4PHI1Z2_L4D4PHI2Z2_SP_L3D4PHI1Z2_L4D4PHI2Z2_wr_en),
.number_out(SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI2Z2_L4D4PHI2Z2_SP_L3D4PHI2Z2_L4D4PHI2Z2;
wire TE_L3D4PHI2Z2_L4D4PHI2Z2_SP_L3D4PHI2Z2_L4D4PHI2Z2_wr_en;
wire [5:0] SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2Z2_L4D4PHI2Z2(
.data_in(TE_L3D4PHI2Z2_L4D4PHI2Z2_SP_L3D4PHI2Z2_L4D4PHI2Z2),
.enable(TE_L3D4PHI2Z2_L4D4PHI2Z2_SP_L3D4PHI2Z2_L4D4PHI2Z2_wr_en),
.number_out(SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI2Z2_L4D4PHI3Z2_SP_L3D4PHI2Z2_L4D4PHI3Z2;
wire TE_L3D4PHI2Z2_L4D4PHI3Z2_SP_L3D4PHI2Z2_L4D4PHI3Z2_wr_en;
wire [5:0] SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2Z2_L4D4PHI3Z2(
.data_in(TE_L3D4PHI2Z2_L4D4PHI3Z2_SP_L3D4PHI2Z2_L4D4PHI3Z2),
.enable(TE_L3D4PHI2Z2_L4D4PHI3Z2_SP_L3D4PHI2Z2_L4D4PHI3Z2_wr_en),
.number_out(SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI3Z2_L4D4PHI3Z2_SP_L3D4PHI3Z2_L4D4PHI3Z2;
wire TE_L3D4PHI3Z2_L4D4PHI3Z2_SP_L3D4PHI3Z2_L4D4PHI3Z2_wr_en;
wire [5:0] SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3Z2_L4D4PHI3Z2(
.data_in(TE_L3D4PHI3Z2_L4D4PHI3Z2_SP_L3D4PHI3Z2_L4D4PHI3Z2),
.enable(TE_L3D4PHI3Z2_L4D4PHI3Z2_SP_L3D4PHI3Z2_L4D4PHI3Z2_wr_en),
.number_out(SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L3D4PHI3Z2_L4D4PHI4Z2_SP_L3D4PHI3Z2_L4D4PHI4Z2;
wire TE_L3D4PHI3Z2_L4D4PHI4Z2_SP_L3D4PHI3Z2_L4D4PHI4Z2_wr_en;
wire [5:0] SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3Z2_L4D4PHI4Z2(
.data_in(TE_L3D4PHI3Z2_L4D4PHI4Z2_SP_L3D4PHI3Z2_L4D4PHI4Z2),
.enable(TE_L3D4PHI3Z2_L4D4PHI4Z2_SP_L3D4PHI3Z2_L4D4PHI4Z2_wr_en),
.number_out(SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L3D4_AS_L3D4n1;
wire VMR_L3D4_AS_L3D4n1_wr_en;
wire [10:0] AS_L3D4n1_TC_L3D4L4D4_read_add;
wire [35:0] AS_L3D4n1_TC_L3D4L4D4;
AllStubs  AS_L3D4n1(
.data_in(VMR_L3D4_AS_L3D4n1),
.enable(VMR_L3D4_AS_L3D4n1_wr_en),
.read_add(AS_L3D4n1_TC_L3D4L4D4_read_add),
.data_out(AS_L3D4n1_TC_L3D4L4D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L4D4_AS_L4D4n2;
wire VMR_L4D4_AS_L4D4n2_wr_en;
wire [10:0] AS_L4D4n2_TC_L3D4L4D4_read_add;
wire [35:0] AS_L4D4n2_TC_L3D4L4D4;
AllStubs  AS_L4D4n2(
.data_in(VMR_L4D4_AS_L4D4n2),
.enable(VMR_L4D4_AS_L4D4n2_wr_en),
.read_add(AS_L4D4n2_TC_L3D4L4D4_read_add),
.data_out(AS_L4D4n2_TC_L3D4L4D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI1Z1_L6D3PHI1Z1_SP_L5D3PHI1Z1_L6D3PHI1Z1;
wire TE_L5D3PHI1Z1_L6D3PHI1Z1_SP_L5D3PHI1Z1_L6D3PHI1Z1_wr_en;
wire [5:0] SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1Z1_L6D3PHI1Z1(
.data_in(TE_L5D3PHI1Z1_L6D3PHI1Z1_SP_L5D3PHI1Z1_L6D3PHI1Z1),
.enable(TE_L5D3PHI1Z1_L6D3PHI1Z1_SP_L5D3PHI1Z1_L6D3PHI1Z1_wr_en),
.number_out(SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI1Z1_L6D3PHI2Z1_SP_L5D3PHI1Z1_L6D3PHI2Z1;
wire TE_L5D3PHI1Z1_L6D3PHI2Z1_SP_L5D3PHI1Z1_L6D3PHI2Z1_wr_en;
wire [5:0] SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1Z1_L6D3PHI2Z1(
.data_in(TE_L5D3PHI1Z1_L6D3PHI2Z1_SP_L5D3PHI1Z1_L6D3PHI2Z1),
.enable(TE_L5D3PHI1Z1_L6D3PHI2Z1_SP_L5D3PHI1Z1_L6D3PHI2Z1_wr_en),
.number_out(SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI2Z1_L6D3PHI2Z1_SP_L5D3PHI2Z1_L6D3PHI2Z1;
wire TE_L5D3PHI2Z1_L6D3PHI2Z1_SP_L5D3PHI2Z1_L6D3PHI2Z1_wr_en;
wire [5:0] SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2Z1_L6D3PHI2Z1(
.data_in(TE_L5D3PHI2Z1_L6D3PHI2Z1_SP_L5D3PHI2Z1_L6D3PHI2Z1),
.enable(TE_L5D3PHI2Z1_L6D3PHI2Z1_SP_L5D3PHI2Z1_L6D3PHI2Z1_wr_en),
.number_out(SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI2Z1_L6D3PHI3Z1_SP_L5D3PHI2Z1_L6D3PHI3Z1;
wire TE_L5D3PHI2Z1_L6D3PHI3Z1_SP_L5D3PHI2Z1_L6D3PHI3Z1_wr_en;
wire [5:0] SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2Z1_L6D3PHI3Z1(
.data_in(TE_L5D3PHI2Z1_L6D3PHI3Z1_SP_L5D3PHI2Z1_L6D3PHI3Z1),
.enable(TE_L5D3PHI2Z1_L6D3PHI3Z1_SP_L5D3PHI2Z1_L6D3PHI3Z1_wr_en),
.number_out(SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI3Z1_L6D3PHI3Z1_SP_L5D3PHI3Z1_L6D3PHI3Z1;
wire TE_L5D3PHI3Z1_L6D3PHI3Z1_SP_L5D3PHI3Z1_L6D3PHI3Z1_wr_en;
wire [5:0] SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3Z1_L6D3PHI3Z1(
.data_in(TE_L5D3PHI3Z1_L6D3PHI3Z1_SP_L5D3PHI3Z1_L6D3PHI3Z1),
.enable(TE_L5D3PHI3Z1_L6D3PHI3Z1_SP_L5D3PHI3Z1_L6D3PHI3Z1_wr_en),
.number_out(SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI3Z1_L6D3PHI4Z1_SP_L5D3PHI3Z1_L6D3PHI4Z1;
wire TE_L5D3PHI3Z1_L6D3PHI4Z1_SP_L5D3PHI3Z1_L6D3PHI4Z1_wr_en;
wire [5:0] SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3Z1_L6D3PHI4Z1(
.data_in(TE_L5D3PHI3Z1_L6D3PHI4Z1_SP_L5D3PHI3Z1_L6D3PHI4Z1),
.enable(TE_L5D3PHI3Z1_L6D3PHI4Z1_SP_L5D3PHI3Z1_L6D3PHI4Z1_wr_en),
.number_out(SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI1Z1_L6D3PHI1Z2_SP_L5D3PHI1Z1_L6D3PHI1Z2;
wire TE_L5D3PHI1Z1_L6D3PHI1Z2_SP_L5D3PHI1Z1_L6D3PHI1Z2_wr_en;
wire [5:0] SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1Z1_L6D3PHI1Z2(
.data_in(TE_L5D3PHI1Z1_L6D3PHI1Z2_SP_L5D3PHI1Z1_L6D3PHI1Z2),
.enable(TE_L5D3PHI1Z1_L6D3PHI1Z2_SP_L5D3PHI1Z1_L6D3PHI1Z2_wr_en),
.number_out(SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI1Z1_L6D3PHI2Z2_SP_L5D3PHI1Z1_L6D3PHI2Z2;
wire TE_L5D3PHI1Z1_L6D3PHI2Z2_SP_L5D3PHI1Z1_L6D3PHI2Z2_wr_en;
wire [5:0] SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1Z1_L6D3PHI2Z2(
.data_in(TE_L5D3PHI1Z1_L6D3PHI2Z2_SP_L5D3PHI1Z1_L6D3PHI2Z2),
.enable(TE_L5D3PHI1Z1_L6D3PHI2Z2_SP_L5D3PHI1Z1_L6D3PHI2Z2_wr_en),
.number_out(SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI2Z1_L6D3PHI2Z2_SP_L5D3PHI2Z1_L6D3PHI2Z2;
wire TE_L5D3PHI2Z1_L6D3PHI2Z2_SP_L5D3PHI2Z1_L6D3PHI2Z2_wr_en;
wire [5:0] SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2Z1_L6D3PHI2Z2(
.data_in(TE_L5D3PHI2Z1_L6D3PHI2Z2_SP_L5D3PHI2Z1_L6D3PHI2Z2),
.enable(TE_L5D3PHI2Z1_L6D3PHI2Z2_SP_L5D3PHI2Z1_L6D3PHI2Z2_wr_en),
.number_out(SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI2Z1_L6D3PHI3Z2_SP_L5D3PHI2Z1_L6D3PHI3Z2;
wire TE_L5D3PHI2Z1_L6D3PHI3Z2_SP_L5D3PHI2Z1_L6D3PHI3Z2_wr_en;
wire [5:0] SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2Z1_L6D3PHI3Z2(
.data_in(TE_L5D3PHI2Z1_L6D3PHI3Z2_SP_L5D3PHI2Z1_L6D3PHI3Z2),
.enable(TE_L5D3PHI2Z1_L6D3PHI3Z2_SP_L5D3PHI2Z1_L6D3PHI3Z2_wr_en),
.number_out(SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI3Z1_L6D3PHI3Z2_SP_L5D3PHI3Z1_L6D3PHI3Z2;
wire TE_L5D3PHI3Z1_L6D3PHI3Z2_SP_L5D3PHI3Z1_L6D3PHI3Z2_wr_en;
wire [5:0] SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3Z1_L6D3PHI3Z2(
.data_in(TE_L5D3PHI3Z1_L6D3PHI3Z2_SP_L5D3PHI3Z1_L6D3PHI3Z2),
.enable(TE_L5D3PHI3Z1_L6D3PHI3Z2_SP_L5D3PHI3Z1_L6D3PHI3Z2_wr_en),
.number_out(SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI3Z1_L6D3PHI4Z2_SP_L5D3PHI3Z1_L6D3PHI4Z2;
wire TE_L5D3PHI3Z1_L6D3PHI4Z2_SP_L5D3PHI3Z1_L6D3PHI4Z2_wr_en;
wire [5:0] SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3Z1_L6D3PHI4Z2(
.data_in(TE_L5D3PHI3Z1_L6D3PHI4Z2_SP_L5D3PHI3Z1_L6D3PHI4Z2),
.enable(TE_L5D3PHI3Z1_L6D3PHI4Z2_SP_L5D3PHI3Z1_L6D3PHI4Z2_wr_en),
.number_out(SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI1Z2_L6D3PHI1Z2_SP_L5D3PHI1Z2_L6D3PHI1Z2;
wire TE_L5D3PHI1Z2_L6D3PHI1Z2_SP_L5D3PHI1Z2_L6D3PHI1Z2_wr_en;
wire [5:0] SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1Z2_L6D3PHI1Z2(
.data_in(TE_L5D3PHI1Z2_L6D3PHI1Z2_SP_L5D3PHI1Z2_L6D3PHI1Z2),
.enable(TE_L5D3PHI1Z2_L6D3PHI1Z2_SP_L5D3PHI1Z2_L6D3PHI1Z2_wr_en),
.number_out(SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI1Z2_L6D3PHI2Z2_SP_L5D3PHI1Z2_L6D3PHI2Z2;
wire TE_L5D3PHI1Z2_L6D3PHI2Z2_SP_L5D3PHI1Z2_L6D3PHI2Z2_wr_en;
wire [5:0] SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1Z2_L6D3PHI2Z2(
.data_in(TE_L5D3PHI1Z2_L6D3PHI2Z2_SP_L5D3PHI1Z2_L6D3PHI2Z2),
.enable(TE_L5D3PHI1Z2_L6D3PHI2Z2_SP_L5D3PHI1Z2_L6D3PHI2Z2_wr_en),
.number_out(SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI2Z2_L6D3PHI2Z2_SP_L5D3PHI2Z2_L6D3PHI2Z2;
wire TE_L5D3PHI2Z2_L6D3PHI2Z2_SP_L5D3PHI2Z2_L6D3PHI2Z2_wr_en;
wire [5:0] SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2Z2_L6D3PHI2Z2(
.data_in(TE_L5D3PHI2Z2_L6D3PHI2Z2_SP_L5D3PHI2Z2_L6D3PHI2Z2),
.enable(TE_L5D3PHI2Z2_L6D3PHI2Z2_SP_L5D3PHI2Z2_L6D3PHI2Z2_wr_en),
.number_out(SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI2Z2_L6D3PHI3Z2_SP_L5D3PHI2Z2_L6D3PHI3Z2;
wire TE_L5D3PHI2Z2_L6D3PHI3Z2_SP_L5D3PHI2Z2_L6D3PHI3Z2_wr_en;
wire [5:0] SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2Z2_L6D3PHI3Z2(
.data_in(TE_L5D3PHI2Z2_L6D3PHI3Z2_SP_L5D3PHI2Z2_L6D3PHI3Z2),
.enable(TE_L5D3PHI2Z2_L6D3PHI3Z2_SP_L5D3PHI2Z2_L6D3PHI3Z2_wr_en),
.number_out(SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI3Z2_L6D3PHI3Z2_SP_L5D3PHI3Z2_L6D3PHI3Z2;
wire TE_L5D3PHI3Z2_L6D3PHI3Z2_SP_L5D3PHI3Z2_L6D3PHI3Z2_wr_en;
wire [5:0] SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3Z2_L6D3PHI3Z2(
.data_in(TE_L5D3PHI3Z2_L6D3PHI3Z2_SP_L5D3PHI3Z2_L6D3PHI3Z2),
.enable(TE_L5D3PHI3Z2_L6D3PHI3Z2_SP_L5D3PHI3Z2_L6D3PHI3Z2_wr_en),
.number_out(SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI3Z2_L6D3PHI4Z2_SP_L5D3PHI3Z2_L6D3PHI4Z2;
wire TE_L5D3PHI3Z2_L6D3PHI4Z2_SP_L5D3PHI3Z2_L6D3PHI4Z2_wr_en;
wire [5:0] SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3Z2_L6D3PHI4Z2(
.data_in(TE_L5D3PHI3Z2_L6D3PHI4Z2_SP_L5D3PHI3Z2_L6D3PHI4Z2),
.enable(TE_L5D3PHI3Z2_L6D3PHI4Z2_SP_L5D3PHI3Z2_L6D3PHI4Z2_wr_en),
.number_out(SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L5D3_AS_L5D3n1;
wire VMR_L5D3_AS_L5D3n1_wr_en;
wire [10:0] AS_L5D3n1_TC_L5D3L6D3_read_add;
wire [35:0] AS_L5D3n1_TC_L5D3L6D3;
AllStubs  AS_L5D3n1(
.data_in(VMR_L5D3_AS_L5D3n1),
.enable(VMR_L5D3_AS_L5D3n1_wr_en),
.read_add(AS_L5D3n1_TC_L5D3L6D3_read_add),
.data_out(AS_L5D3n1_TC_L5D3L6D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L6D3_AS_L6D3n1;
wire VMR_L6D3_AS_L6D3n1_wr_en;
wire [10:0] AS_L6D3n1_TC_L5D3L6D3_read_add;
wire [35:0] AS_L6D3n1_TC_L5D3L6D3;
AllStubs  AS_L6D3n1(
.data_in(VMR_L6D3_AS_L6D3n1),
.enable(VMR_L6D3_AS_L6D3n1_wr_en),
.read_add(AS_L6D3n1_TC_L5D3L6D3_read_add),
.data_out(AS_L6D3n1_TC_L5D3L6D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI1Z2_L6D4PHI1Z1_SP_L5D3PHI1Z2_L6D4PHI1Z1;
wire TE_L5D3PHI1Z2_L6D4PHI1Z1_SP_L5D3PHI1Z2_L6D4PHI1Z1_wr_en;
wire [5:0] SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI1Z2_L6D4PHI1Z1(
.data_in(TE_L5D3PHI1Z2_L6D4PHI1Z1_SP_L5D3PHI1Z2_L6D4PHI1Z1),
.enable(TE_L5D3PHI1Z2_L6D4PHI1Z1_SP_L5D3PHI1Z2_L6D4PHI1Z1_wr_en),
.number_out(SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI1Z2_L6D4PHI2Z1_SP_L5D3PHI1Z2_L6D4PHI2Z1;
wire TE_L5D3PHI1Z2_L6D4PHI2Z1_SP_L5D3PHI1Z2_L6D4PHI2Z1_wr_en;
wire [5:0] SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI1Z2_L6D4PHI2Z1(
.data_in(TE_L5D3PHI1Z2_L6D4PHI2Z1_SP_L5D3PHI1Z2_L6D4PHI2Z1),
.enable(TE_L5D3PHI1Z2_L6D4PHI2Z1_SP_L5D3PHI1Z2_L6D4PHI2Z1_wr_en),
.number_out(SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI2Z2_L6D4PHI2Z1_SP_L5D3PHI2Z2_L6D4PHI2Z1;
wire TE_L5D3PHI2Z2_L6D4PHI2Z1_SP_L5D3PHI2Z2_L6D4PHI2Z1_wr_en;
wire [5:0] SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI2Z2_L6D4PHI2Z1(
.data_in(TE_L5D3PHI2Z2_L6D4PHI2Z1_SP_L5D3PHI2Z2_L6D4PHI2Z1),
.enable(TE_L5D3PHI2Z2_L6D4PHI2Z1_SP_L5D3PHI2Z2_L6D4PHI2Z1_wr_en),
.number_out(SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI2Z2_L6D4PHI3Z1_SP_L5D3PHI2Z2_L6D4PHI3Z1;
wire TE_L5D3PHI2Z2_L6D4PHI3Z1_SP_L5D3PHI2Z2_L6D4PHI3Z1_wr_en;
wire [5:0] SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI2Z2_L6D4PHI3Z1(
.data_in(TE_L5D3PHI2Z2_L6D4PHI3Z1_SP_L5D3PHI2Z2_L6D4PHI3Z1),
.enable(TE_L5D3PHI2Z2_L6D4PHI3Z1_SP_L5D3PHI2Z2_L6D4PHI3Z1_wr_en),
.number_out(SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI3Z2_L6D4PHI3Z1_SP_L5D3PHI3Z2_L6D4PHI3Z1;
wire TE_L5D3PHI3Z2_L6D4PHI3Z1_SP_L5D3PHI3Z2_L6D4PHI3Z1_wr_en;
wire [5:0] SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI3Z2_L6D4PHI3Z1(
.data_in(TE_L5D3PHI3Z2_L6D4PHI3Z1_SP_L5D3PHI3Z2_L6D4PHI3Z1),
.enable(TE_L5D3PHI3Z2_L6D4PHI3Z1_SP_L5D3PHI3Z2_L6D4PHI3Z1_wr_en),
.number_out(SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D3PHI3Z2_L6D4PHI4Z1_SP_L5D3PHI3Z2_L6D4PHI4Z1;
wire TE_L5D3PHI3Z2_L6D4PHI4Z1_SP_L5D3PHI3Z2_L6D4PHI4Z1_wr_en;
wire [5:0] SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI3Z2_L6D4PHI4Z1(
.data_in(TE_L5D3PHI3Z2_L6D4PHI4Z1_SP_L5D3PHI3Z2_L6D4PHI4Z1),
.enable(TE_L5D3PHI3Z2_L6D4PHI4Z1_SP_L5D3PHI3Z2_L6D4PHI4Z1_wr_en),
.number_out(SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L5D3_AS_L5D3n2;
wire VMR_L5D3_AS_L5D3n2_wr_en;
wire [10:0] AS_L5D3n2_TC_L5D3L6D4_read_add;
wire [35:0] AS_L5D3n2_TC_L5D3L6D4;
AllStubs  AS_L5D3n2(
.data_in(VMR_L5D3_AS_L5D3n2),
.enable(VMR_L5D3_AS_L5D3n2_wr_en),
.read_add(AS_L5D3n2_TC_L5D3L6D4_read_add),
.data_out(AS_L5D3n2_TC_L5D3L6D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L6D4_AS_L6D4n1;
wire VMR_L6D4_AS_L6D4n1_wr_en;
wire [10:0] AS_L6D4n1_TC_L5D3L6D4_read_add;
wire [35:0] AS_L6D4n1_TC_L5D3L6D4;
AllStubs  AS_L6D4n1(
.data_in(VMR_L6D4_AS_L6D4n1),
.enable(VMR_L6D4_AS_L6D4n1_wr_en),
.read_add(AS_L6D4n1_TC_L5D3L6D4_read_add),
.data_out(AS_L6D4n1_TC_L5D3L6D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI1Z1_L6D4PHI1Z1_SP_L5D4PHI1Z1_L6D4PHI1Z1;
wire TE_L5D4PHI1Z1_L6D4PHI1Z1_SP_L5D4PHI1Z1_L6D4PHI1Z1_wr_en;
wire [5:0] SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1Z1_L6D4PHI1Z1(
.data_in(TE_L5D4PHI1Z1_L6D4PHI1Z1_SP_L5D4PHI1Z1_L6D4PHI1Z1),
.enable(TE_L5D4PHI1Z1_L6D4PHI1Z1_SP_L5D4PHI1Z1_L6D4PHI1Z1_wr_en),
.number_out(SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI1Z1_L6D4PHI2Z1_SP_L5D4PHI1Z1_L6D4PHI2Z1;
wire TE_L5D4PHI1Z1_L6D4PHI2Z1_SP_L5D4PHI1Z1_L6D4PHI2Z1_wr_en;
wire [5:0] SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1Z1_L6D4PHI2Z1(
.data_in(TE_L5D4PHI1Z1_L6D4PHI2Z1_SP_L5D4PHI1Z1_L6D4PHI2Z1),
.enable(TE_L5D4PHI1Z1_L6D4PHI2Z1_SP_L5D4PHI1Z1_L6D4PHI2Z1_wr_en),
.number_out(SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI2Z1_L6D4PHI2Z1_SP_L5D4PHI2Z1_L6D4PHI2Z1;
wire TE_L5D4PHI2Z1_L6D4PHI2Z1_SP_L5D4PHI2Z1_L6D4PHI2Z1_wr_en;
wire [5:0] SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2Z1_L6D4PHI2Z1(
.data_in(TE_L5D4PHI2Z1_L6D4PHI2Z1_SP_L5D4PHI2Z1_L6D4PHI2Z1),
.enable(TE_L5D4PHI2Z1_L6D4PHI2Z1_SP_L5D4PHI2Z1_L6D4PHI2Z1_wr_en),
.number_out(SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI2Z1_L6D4PHI3Z1_SP_L5D4PHI2Z1_L6D4PHI3Z1;
wire TE_L5D4PHI2Z1_L6D4PHI3Z1_SP_L5D4PHI2Z1_L6D4PHI3Z1_wr_en;
wire [5:0] SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2Z1_L6D4PHI3Z1(
.data_in(TE_L5D4PHI2Z1_L6D4PHI3Z1_SP_L5D4PHI2Z1_L6D4PHI3Z1),
.enable(TE_L5D4PHI2Z1_L6D4PHI3Z1_SP_L5D4PHI2Z1_L6D4PHI3Z1_wr_en),
.number_out(SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI3Z1_L6D4PHI3Z1_SP_L5D4PHI3Z1_L6D4PHI3Z1;
wire TE_L5D4PHI3Z1_L6D4PHI3Z1_SP_L5D4PHI3Z1_L6D4PHI3Z1_wr_en;
wire [5:0] SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3Z1_L6D4PHI3Z1(
.data_in(TE_L5D4PHI3Z1_L6D4PHI3Z1_SP_L5D4PHI3Z1_L6D4PHI3Z1),
.enable(TE_L5D4PHI3Z1_L6D4PHI3Z1_SP_L5D4PHI3Z1_L6D4PHI3Z1_wr_en),
.number_out(SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI3Z1_L6D4PHI4Z1_SP_L5D4PHI3Z1_L6D4PHI4Z1;
wire TE_L5D4PHI3Z1_L6D4PHI4Z1_SP_L5D4PHI3Z1_L6D4PHI4Z1_wr_en;
wire [5:0] SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3Z1_L6D4PHI4Z1(
.data_in(TE_L5D4PHI3Z1_L6D4PHI4Z1_SP_L5D4PHI3Z1_L6D4PHI4Z1),
.enable(TE_L5D4PHI3Z1_L6D4PHI4Z1_SP_L5D4PHI3Z1_L6D4PHI4Z1_wr_en),
.number_out(SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI1Z1_L6D4PHI1Z2_SP_L5D4PHI1Z1_L6D4PHI1Z2;
wire TE_L5D4PHI1Z1_L6D4PHI1Z2_SP_L5D4PHI1Z1_L6D4PHI1Z2_wr_en;
wire [5:0] SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1Z1_L6D4PHI1Z2(
.data_in(TE_L5D4PHI1Z1_L6D4PHI1Z2_SP_L5D4PHI1Z1_L6D4PHI1Z2),
.enable(TE_L5D4PHI1Z1_L6D4PHI1Z2_SP_L5D4PHI1Z1_L6D4PHI1Z2_wr_en),
.number_out(SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI1Z1_L6D4PHI2Z2_SP_L5D4PHI1Z1_L6D4PHI2Z2;
wire TE_L5D4PHI1Z1_L6D4PHI2Z2_SP_L5D4PHI1Z1_L6D4PHI2Z2_wr_en;
wire [5:0] SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1Z1_L6D4PHI2Z2(
.data_in(TE_L5D4PHI1Z1_L6D4PHI2Z2_SP_L5D4PHI1Z1_L6D4PHI2Z2),
.enable(TE_L5D4PHI1Z1_L6D4PHI2Z2_SP_L5D4PHI1Z1_L6D4PHI2Z2_wr_en),
.number_out(SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI2Z1_L6D4PHI2Z2_SP_L5D4PHI2Z1_L6D4PHI2Z2;
wire TE_L5D4PHI2Z1_L6D4PHI2Z2_SP_L5D4PHI2Z1_L6D4PHI2Z2_wr_en;
wire [5:0] SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2Z1_L6D4PHI2Z2(
.data_in(TE_L5D4PHI2Z1_L6D4PHI2Z2_SP_L5D4PHI2Z1_L6D4PHI2Z2),
.enable(TE_L5D4PHI2Z1_L6D4PHI2Z2_SP_L5D4PHI2Z1_L6D4PHI2Z2_wr_en),
.number_out(SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI2Z1_L6D4PHI3Z2_SP_L5D4PHI2Z1_L6D4PHI3Z2;
wire TE_L5D4PHI2Z1_L6D4PHI3Z2_SP_L5D4PHI2Z1_L6D4PHI3Z2_wr_en;
wire [5:0] SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2Z1_L6D4PHI3Z2(
.data_in(TE_L5D4PHI2Z1_L6D4PHI3Z2_SP_L5D4PHI2Z1_L6D4PHI3Z2),
.enable(TE_L5D4PHI2Z1_L6D4PHI3Z2_SP_L5D4PHI2Z1_L6D4PHI3Z2_wr_en),
.number_out(SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI3Z1_L6D4PHI3Z2_SP_L5D4PHI3Z1_L6D4PHI3Z2;
wire TE_L5D4PHI3Z1_L6D4PHI3Z2_SP_L5D4PHI3Z1_L6D4PHI3Z2_wr_en;
wire [5:0] SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3Z1_L6D4PHI3Z2(
.data_in(TE_L5D4PHI3Z1_L6D4PHI3Z2_SP_L5D4PHI3Z1_L6D4PHI3Z2),
.enable(TE_L5D4PHI3Z1_L6D4PHI3Z2_SP_L5D4PHI3Z1_L6D4PHI3Z2_wr_en),
.number_out(SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI3Z1_L6D4PHI4Z2_SP_L5D4PHI3Z1_L6D4PHI4Z2;
wire TE_L5D4PHI3Z1_L6D4PHI4Z2_SP_L5D4PHI3Z1_L6D4PHI4Z2_wr_en;
wire [5:0] SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3Z1_L6D4PHI4Z2(
.data_in(TE_L5D4PHI3Z1_L6D4PHI4Z2_SP_L5D4PHI3Z1_L6D4PHI4Z2),
.enable(TE_L5D4PHI3Z1_L6D4PHI4Z2_SP_L5D4PHI3Z1_L6D4PHI4Z2_wr_en),
.number_out(SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI1Z2_L6D4PHI1Z2_SP_L5D4PHI1Z2_L6D4PHI1Z2;
wire TE_L5D4PHI1Z2_L6D4PHI1Z2_SP_L5D4PHI1Z2_L6D4PHI1Z2_wr_en;
wire [5:0] SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1Z2_L6D4PHI1Z2(
.data_in(TE_L5D4PHI1Z2_L6D4PHI1Z2_SP_L5D4PHI1Z2_L6D4PHI1Z2),
.enable(TE_L5D4PHI1Z2_L6D4PHI1Z2_SP_L5D4PHI1Z2_L6D4PHI1Z2_wr_en),
.number_out(SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI1Z2_L6D4PHI2Z2_SP_L5D4PHI1Z2_L6D4PHI2Z2;
wire TE_L5D4PHI1Z2_L6D4PHI2Z2_SP_L5D4PHI1Z2_L6D4PHI2Z2_wr_en;
wire [5:0] SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1Z2_L6D4PHI2Z2(
.data_in(TE_L5D4PHI1Z2_L6D4PHI2Z2_SP_L5D4PHI1Z2_L6D4PHI2Z2),
.enable(TE_L5D4PHI1Z2_L6D4PHI2Z2_SP_L5D4PHI1Z2_L6D4PHI2Z2_wr_en),
.number_out(SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI2Z2_L6D4PHI2Z2_SP_L5D4PHI2Z2_L6D4PHI2Z2;
wire TE_L5D4PHI2Z2_L6D4PHI2Z2_SP_L5D4PHI2Z2_L6D4PHI2Z2_wr_en;
wire [5:0] SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2Z2_L6D4PHI2Z2(
.data_in(TE_L5D4PHI2Z2_L6D4PHI2Z2_SP_L5D4PHI2Z2_L6D4PHI2Z2),
.enable(TE_L5D4PHI2Z2_L6D4PHI2Z2_SP_L5D4PHI2Z2_L6D4PHI2Z2_wr_en),
.number_out(SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI2Z2_L6D4PHI3Z2_SP_L5D4PHI2Z2_L6D4PHI3Z2;
wire TE_L5D4PHI2Z2_L6D4PHI3Z2_SP_L5D4PHI2Z2_L6D4PHI3Z2_wr_en;
wire [5:0] SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2Z2_L6D4PHI3Z2(
.data_in(TE_L5D4PHI2Z2_L6D4PHI3Z2_SP_L5D4PHI2Z2_L6D4PHI3Z2),
.enable(TE_L5D4PHI2Z2_L6D4PHI3Z2_SP_L5D4PHI2Z2_L6D4PHI3Z2_wr_en),
.number_out(SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI3Z2_L6D4PHI3Z2_SP_L5D4PHI3Z2_L6D4PHI3Z2;
wire TE_L5D4PHI3Z2_L6D4PHI3Z2_SP_L5D4PHI3Z2_L6D4PHI3Z2_wr_en;
wire [5:0] SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3Z2_L6D4PHI3Z2(
.data_in(TE_L5D4PHI3Z2_L6D4PHI3Z2_SP_L5D4PHI3Z2_L6D4PHI3Z2),
.enable(TE_L5D4PHI3Z2_L6D4PHI3Z2_SP_L5D4PHI3Z2_L6D4PHI3Z2_wr_en),
.number_out(SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] TE_L5D4PHI3Z2_L6D4PHI4Z2_SP_L5D4PHI3Z2_L6D4PHI4Z2;
wire TE_L5D4PHI3Z2_L6D4PHI4Z2_SP_L5D4PHI3Z2_L6D4PHI4Z2_wr_en;
wire [5:0] SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3Z2_L6D4PHI4Z2(
.data_in(TE_L5D4PHI3Z2_L6D4PHI4Z2_SP_L5D4PHI3Z2_L6D4PHI4Z2),
.enable(TE_L5D4PHI3Z2_L6D4PHI4Z2_SP_L5D4PHI3Z2_L6D4PHI4Z2_wr_en),
.number_out(SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4),
.start(start4_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L5D4_AS_L5D4n1;
wire VMR_L5D4_AS_L5D4n1_wr_en;
wire [10:0] AS_L5D4n1_TC_L5D4L6D4_read_add;
wire [35:0] AS_L5D4n1_TC_L5D4L6D4;
AllStubs  AS_L5D4n1(
.data_in(VMR_L5D4_AS_L5D4n1),
.enable(VMR_L5D4_AS_L5D4n1_wr_en),
.read_add(AS_L5D4n1_TC_L5D4L6D4_read_add),
.data_out(AS_L5D4n1_TC_L5D4L6D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L6D4_AS_L6D4n2;
wire VMR_L6D4_AS_L6D4n2_wr_en;
wire [10:0] AS_L6D4n2_TC_L5D4L6D4_read_add;
wire [35:0] AS_L6D4n2_TC_L5D4L6D4;
AllStubs  AS_L6D4n2(
.data_in(VMR_L6D4_AS_L6D4n2),
.enable(VMR_L6D4_AS_L6D4n2_wr_en),
.read_add(AS_L6D4n2_TC_L5D4L6D4_read_add),
.data_out(AS_L6D4n2_TC_L5D4L6D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3;
wire TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D3L2D3_L3(
.data_in(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3),
.enable(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus),
.start(startproj5_0),
.done(done4_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4;
wire TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D3L2D3_L4(
.data_in(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4),
.enable(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5;
wire TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D3L2D3_L5(
.data_in(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5),
.enable(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6;
wire TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D3L2D3_L6(
.data_in(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6),
.enable(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3;
wire TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D3L2D4_L3(
.data_in(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3),
.enable(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4;
wire TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D3L2D4_L4(
.data_in(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4),
.enable(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L5;
wire TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D3L2D4_L5(
.data_in(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L5),
.enable(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L5_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L6;
wire TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D3L2D4_L6(
.data_in(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L6),
.enable(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L6_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3;
wire TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D4L2D4_L3(
.data_in(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3),
.enable(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3_wr_en),
.number_out(TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L4;
wire TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D4L2D4_L4(
.data_in(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L4),
.enable(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L4_wr_en),
.number_out(TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L5;
wire TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D4L2D4_L5(
.data_in(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L5),
.enable(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L5_wr_en),
.number_out(TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L6;
wire TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus;
TrackletProjections  TPROJ_ToPlus_L1D4L2D4_L6(
.data_in(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L6),
.enable(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L6_wr_en),
.number_out(TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus_number),
.read_add(TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1;
wire TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D3L4D3_L1(
.data_in(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1),
.enable(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2;
wire TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D3L4D3_L2(
.data_in(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2),
.enable(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5;
wire TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D3L4D3_L5(
.data_in(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5),
.enable(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6;
wire TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D3L4D3_L6(
.data_in(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6),
.enable(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1;
wire TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D3L4D4_L1(
.data_in(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1),
.enable(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2;
wire TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D3L4D4_L2(
.data_in(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2),
.enable(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5;
wire TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D3L4D4_L5(
.data_in(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5),
.enable(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6;
wire TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D3L4D4_L6(
.data_in(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6),
.enable(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1;
wire TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D4L4D4_L1(
.data_in(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1),
.enable(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1_wr_en),
.number_out(TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2;
wire TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D4L4D4_L2(
.data_in(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2),
.enable(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2_wr_en),
.number_out(TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5;
wire TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D4L4D4_L5(
.data_in(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5),
.enable(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5_wr_en),
.number_out(TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6;
wire TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus;
TrackletProjections  TPROJ_ToPlus_L3D4L4D4_L6(
.data_in(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6),
.enable(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6_wr_en),
.number_out(TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus_number),
.read_add(TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1;
wire TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D3L6D3_L1(
.data_in(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1),
.enable(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2;
wire TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D3L6D3_L2(
.data_in(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2),
.enable(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3;
wire TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D3L6D3_L3(
.data_in(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3),
.enable(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4;
wire TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D3L6D3_L4(
.data_in(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4),
.enable(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1;
wire TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D3L6D4_L1(
.data_in(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1),
.enable(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2;
wire TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D3L6D4_L2(
.data_in(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2),
.enable(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3;
wire TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D3L6D4_L3(
.data_in(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3),
.enable(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4;
wire TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D3L6D4_L4(
.data_in(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4),
.enable(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1;
wire TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D4L6D4_L1(
.data_in(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1),
.enable(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1_wr_en),
.number_out(TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2;
wire TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D4L6D4_L2(
.data_in(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2),
.enable(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2_wr_en),
.number_out(TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3;
wire TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D4L6D4_L3(
.data_in(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3),
.enable(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3_wr_en),
.number_out(TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4;
wire TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus;
TrackletProjections  TPROJ_ToPlus_L5D4L6D4_L4(
.data_in(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4),
.enable(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4_wr_en),
.number_out(TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus_number),
.read_add(TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3;
wire TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D3L2D3_L3(
.data_in(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3),
.enable(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4;
wire TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D3L2D3_L4(
.data_in(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4),
.enable(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5;
wire TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D3L2D3_L5(
.data_in(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5),
.enable(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6;
wire TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D3L2D3_L6(
.data_in(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6),
.enable(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3;
wire TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D3L2D4_L3(
.data_in(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3),
.enable(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4;
wire TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D3L2D4_L4(
.data_in(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4),
.enable(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L5;
wire TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D3L2D4_L5(
.data_in(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L5),
.enable(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L5_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L6;
wire TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D3L2D4_L6(
.data_in(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L6),
.enable(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L6_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3;
wire TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D4L2D4_L3(
.data_in(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3),
.enable(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3_wr_en),
.number_out(TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L4;
wire TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D4L2D4_L4(
.data_in(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L4),
.enable(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L4_wr_en),
.number_out(TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L5;
wire TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D4L2D4_L5(
.data_in(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L5),
.enable(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L5_wr_en),
.number_out(TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L6;
wire TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus;
TrackletProjections  TPROJ_ToMinus_L1D4L2D4_L6(
.data_in(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L6),
.enable(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L6_wr_en),
.number_out(TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus_number),
.read_add(TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1;
wire TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D3L4D3_L1(
.data_in(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1),
.enable(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2;
wire TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D3L4D3_L2(
.data_in(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2),
.enable(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5;
wire TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D3L4D3_L5(
.data_in(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5),
.enable(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6;
wire TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D3L4D3_L6(
.data_in(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6),
.enable(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1;
wire TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D3L4D4_L1(
.data_in(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1),
.enable(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2;
wire TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D3L4D4_L2(
.data_in(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2),
.enable(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5;
wire TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D3L4D4_L5(
.data_in(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5),
.enable(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6;
wire TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D3L4D4_L6(
.data_in(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6),
.enable(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1;
wire TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D4L4D4_L1(
.data_in(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1),
.enable(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1_wr_en),
.number_out(TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2;
wire TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D4L4D4_L2(
.data_in(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2),
.enable(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2_wr_en),
.number_out(TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5;
wire TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D4L4D4_L5(
.data_in(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5),
.enable(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5_wr_en),
.number_out(TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6;
wire TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus;
TrackletProjections  TPROJ_ToMinus_L3D4L4D4_L6(
.data_in(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6),
.enable(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6_wr_en),
.number_out(TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus_number),
.read_add(TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1;
wire TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D3L6D3_L1(
.data_in(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1),
.enable(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2;
wire TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D3L6D3_L2(
.data_in(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2),
.enable(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3;
wire TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D3L6D3_L3(
.data_in(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3),
.enable(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4;
wire TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D3L6D3_L4(
.data_in(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4),
.enable(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1;
wire TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D3L6D4_L1(
.data_in(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1),
.enable(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2;
wire TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D3L6D4_L2(
.data_in(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2),
.enable(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3;
wire TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D3L6D4_L3(
.data_in(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3),
.enable(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4;
wire TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D3L6D4_L4(
.data_in(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4),
.enable(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1;
wire TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D4L6D4_L1(
.data_in(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1),
.enable(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1_wr_en),
.number_out(TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2;
wire TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D4L6D4_L2(
.data_in(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2),
.enable(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2_wr_en),
.number_out(TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3;
wire TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D4L6D4_L3(
.data_in(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3),
.enable(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3_wr_en),
.number_out(TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4;
wire TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus;
TrackletProjections  TPROJ_ToMinus_L5D4L6D4_L4(
.data_in(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4),
.enable(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4_wr_en),
.number_out(TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus_number),
.read_add(TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Plus_TPROJ_FromPlus_L1D3_L3L4;
wire PT_L3L4_Plus_TPROJ_FromPlus_L1D3_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4;
TrackletProjections  TPROJ_FromPlus_L1D3_L3L4(
.data_in(PT_L3L4_Plus_TPROJ_FromPlus_L1D3_L3L4),
.enable(PT_L3L4_Plus_TPROJ_FromPlus_L1D3_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_number),
.read_add(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4),
.start(start6_0),
.done(done5_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Minus_TPROJ_FromMinus_L1D3_L3L4;
wire PT_L3L4_Minus_TPROJ_FromMinus_L1D3_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4;
TrackletProjections  TPROJ_FromMinus_L1D3_L3L4(
.data_in(PT_L3L4_Minus_TPROJ_FromMinus_L1D3_L3L4),
.enable(PT_L3L4_Minus_TPROJ_FromMinus_L1D3_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_number),
.read_add(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L1D3(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3_wr_en),
.number_out(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L1D3(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3_wr_en),
.number_out(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L1D3(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3_wr_en),
.number_out(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Plus_TPROJ_FromPlus_L1D4_L3L4;
wire PT_L3L4_Plus_TPROJ_FromPlus_L1D4_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_number;
wire [9:0] TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4;
TrackletProjections  TPROJ_FromPlus_L1D4_L3L4(
.data_in(PT_L3L4_Plus_TPROJ_FromPlus_L1D4_L3L4),
.enable(PT_L3L4_Plus_TPROJ_FromPlus_L1D4_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_number),
.read_add(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_read_add),
.data_out(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Minus_TPROJ_FromMinus_L1D4_L3L4;
wire PT_L3L4_Minus_TPROJ_FromMinus_L1D4_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_number;
wire [9:0] TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4;
TrackletProjections  TPROJ_FromMinus_L1D4_L3L4(
.data_in(PT_L3L4_Minus_TPROJ_FromMinus_L1D4_L3L4),
.enable(PT_L3L4_Minus_TPROJ_FromMinus_L1D4_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_number),
.read_add(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_read_add),
.data_out(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D4;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D4_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L1D4(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D4),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D4_wr_en),
.number_out(TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D4;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D4_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L1D4(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D4),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D4_wr_en),
.number_out(TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D4;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D4_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L1D4(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D4),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D4_wr_en),
.number_out(TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Plus_TPROJ_FromPlus_L2D3_L3L4;
wire PT_L3L4_Plus_TPROJ_FromPlus_L2D3_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4;
TrackletProjections  TPROJ_FromPlus_L2D3_L3L4(
.data_in(PT_L3L4_Plus_TPROJ_FromPlus_L2D3_L3L4),
.enable(PT_L3L4_Plus_TPROJ_FromPlus_L2D3_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_number),
.read_add(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Minus_TPROJ_FromMinus_L2D3_L3L4;
wire PT_L3L4_Minus_TPROJ_FromMinus_L2D3_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4;
TrackletProjections  TPROJ_FromMinus_L2D3_L3L4(
.data_in(PT_L3L4_Minus_TPROJ_FromMinus_L2D3_L3L4),
.enable(PT_L3L4_Minus_TPROJ_FromMinus_L2D3_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_number),
.read_add(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L2D3(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3_wr_en),
.number_out(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L2D3(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3_wr_en),
.number_out(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L2D3(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3_wr_en),
.number_out(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Plus_TPROJ_FromPlus_L2D4_L3L4;
wire PT_L3L4_Plus_TPROJ_FromPlus_L2D4_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_number;
wire [9:0] TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4;
TrackletProjections  TPROJ_FromPlus_L2D4_L3L4(
.data_in(PT_L3L4_Plus_TPROJ_FromPlus_L2D4_L3L4),
.enable(PT_L3L4_Plus_TPROJ_FromPlus_L2D4_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_number),
.read_add(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_read_add),
.data_out(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Minus_TPROJ_FromMinus_L2D4_L3L4;
wire PT_L3L4_Minus_TPROJ_FromMinus_L2D4_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_number;
wire [9:0] TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4;
TrackletProjections  TPROJ_FromMinus_L2D4_L3L4(
.data_in(PT_L3L4_Minus_TPROJ_FromMinus_L2D4_L3L4),
.enable(PT_L3L4_Minus_TPROJ_FromMinus_L2D4_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_number),
.read_add(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_read_add),
.data_out(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D4;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D4_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L2D4(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D4),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D4_wr_en),
.number_out(TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D4;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D4_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L2D4(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D4),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D4_wr_en),
.number_out(TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L2D4(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4_wr_en),
.number_out(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Plus_TPROJ_FromPlus_L5D3_L3L4;
wire PT_L3L4_Plus_TPROJ_FromPlus_L5D3_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_number;
wire [9:0] TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4;
TrackletProjections  TPROJ_FromPlus_L5D3_L3L4(
.data_in(PT_L3L4_Plus_TPROJ_FromPlus_L5D3_L3L4),
.enable(PT_L3L4_Plus_TPROJ_FromPlus_L5D3_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_number),
.read_add(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_read_add),
.data_out(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Minus_TPROJ_FromMinus_L5D3_L3L4;
wire PT_L3L4_Minus_TPROJ_FromMinus_L5D3_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_number;
wire [9:0] TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4;
TrackletProjections  TPROJ_FromMinus_L5D3_L3L4(
.data_in(PT_L3L4_Minus_TPROJ_FromMinus_L5D3_L3L4),
.enable(PT_L3L4_Minus_TPROJ_FromMinus_L5D3_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_number),
.read_add(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_read_add),
.data_out(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L5D3(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3_wr_en),
.number_out(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D3;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D3_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L5D3(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D3),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D3_wr_en),
.number_out(TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D3;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D3_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L5D3(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D3),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D3_wr_en),
.number_out(TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Plus_TPROJ_FromPlus_L5D4_L3L4;
wire PT_L3L4_Plus_TPROJ_FromPlus_L5D4_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4;
TrackletProjections  TPROJ_FromPlus_L5D4_L3L4(
.data_in(PT_L3L4_Plus_TPROJ_FromPlus_L5D4_L3L4),
.enable(PT_L3L4_Plus_TPROJ_FromPlus_L5D4_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_number),
.read_add(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Minus_TPROJ_FromMinus_L5D4_L3L4;
wire PT_L3L4_Minus_TPROJ_FromMinus_L5D4_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4;
TrackletProjections  TPROJ_FromMinus_L5D4_L3L4(
.data_in(PT_L3L4_Minus_TPROJ_FromMinus_L5D4_L3L4),
.enable(PT_L3L4_Minus_TPROJ_FromMinus_L5D4_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_number),
.read_add(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L5D4(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4_wr_en),
.number_out(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L5D4(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4_wr_en),
.number_out(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L5D4(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4_wr_en),
.number_out(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Plus_TPROJ_FromPlus_L6D3_L3L4;
wire PT_L3L4_Plus_TPROJ_FromPlus_L6D3_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_number;
wire [9:0] TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4;
TrackletProjections  TPROJ_FromPlus_L6D3_L3L4(
.data_in(PT_L3L4_Plus_TPROJ_FromPlus_L6D3_L3L4),
.enable(PT_L3L4_Plus_TPROJ_FromPlus_L6D3_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_number),
.read_add(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_read_add),
.data_out(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Minus_TPROJ_FromMinus_L6D3_L3L4;
wire PT_L3L4_Minus_TPROJ_FromMinus_L6D3_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_number;
wire [9:0] TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4;
TrackletProjections  TPROJ_FromMinus_L6D3_L3L4(
.data_in(PT_L3L4_Minus_TPROJ_FromMinus_L6D3_L3L4),
.enable(PT_L3L4_Minus_TPROJ_FromMinus_L6D3_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_number),
.read_add(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_read_add),
.data_out(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L6D3(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3_wr_en),
.number_out(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D3;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D3_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L6D3(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D3),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D3_wr_en),
.number_out(TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D3;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D3_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L6D3(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D3),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D3_wr_en),
.number_out(TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Plus_TPROJ_FromPlus_L6D4_L3L4;
wire PT_L3L4_Plus_TPROJ_FromPlus_L6D4_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4;
TrackletProjections  TPROJ_FromPlus_L6D4_L3L4(
.data_in(PT_L3L4_Plus_TPROJ_FromPlus_L6D4_L3L4),
.enable(PT_L3L4_Plus_TPROJ_FromPlus_L6D4_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_number),
.read_add(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L3L4_Minus_TPROJ_FromMinus_L6D4_L3L4;
wire PT_L3L4_Minus_TPROJ_FromMinus_L6D4_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4;
TrackletProjections  TPROJ_FromMinus_L6D4_L3L4(
.data_in(PT_L3L4_Minus_TPROJ_FromMinus_L6D4_L3L4),
.enable(PT_L3L4_Minus_TPROJ_FromMinus_L6D4_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_number),
.read_add(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L6D4(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4_wr_en),
.number_out(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L6D4(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4_wr_en),
.number_out(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L6D4(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4_wr_en),
.number_out(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Plus_TPROJ_FromPlus_L3D3_L1L2;
wire PT_L1L2_Plus_TPROJ_FromPlus_L3D3_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_number;
wire [9:0] TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2;
TrackletProjections  TPROJ_FromPlus_L3D3_L1L2(
.data_in(PT_L1L2_Plus_TPROJ_FromPlus_L3D3_L1L2),
.enable(PT_L1L2_Plus_TPROJ_FromPlus_L3D3_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_number),
.read_add(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_read_add),
.data_out(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Minus_TPROJ_FromMinus_L3D3_L1L2;
wire PT_L1L2_Minus_TPROJ_FromMinus_L3D3_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_number;
wire [9:0] TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2;
TrackletProjections  TPROJ_FromMinus_L3D3_L1L2(
.data_in(PT_L1L2_Minus_TPROJ_FromMinus_L3D3_L1L2),
.enable(PT_L1L2_Minus_TPROJ_FromMinus_L3D3_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_number),
.read_add(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_read_add),
.data_out(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L3D3(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3_wr_en),
.number_out(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D3;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D3_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L3D3(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D3),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D3_wr_en),
.number_out(TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D3;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D3_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L3D3(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D3),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D3_wr_en),
.number_out(TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Plus_TPROJ_FromPlus_L3D4_L1L2;
wire PT_L1L2_Plus_TPROJ_FromPlus_L3D4_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2;
TrackletProjections  TPROJ_FromPlus_L3D4_L1L2(
.data_in(PT_L1L2_Plus_TPROJ_FromPlus_L3D4_L1L2),
.enable(PT_L1L2_Plus_TPROJ_FromPlus_L3D4_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_number),
.read_add(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Minus_TPROJ_FromMinus_L3D4_L1L2;
wire PT_L1L2_Minus_TPROJ_FromMinus_L3D4_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2;
TrackletProjections  TPROJ_FromMinus_L3D4_L1L2(
.data_in(PT_L1L2_Minus_TPROJ_FromMinus_L3D4_L1L2),
.enable(PT_L1L2_Minus_TPROJ_FromMinus_L3D4_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_number),
.read_add(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L3D4(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4_wr_en),
.number_out(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L3D4(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4_wr_en),
.number_out(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L3D4(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4_wr_en),
.number_out(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Plus_TPROJ_FromPlus_L4D3_L1L2;
wire PT_L1L2_Plus_TPROJ_FromPlus_L4D3_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_number;
wire [9:0] TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2;
TrackletProjections  TPROJ_FromPlus_L4D3_L1L2(
.data_in(PT_L1L2_Plus_TPROJ_FromPlus_L4D3_L1L2),
.enable(PT_L1L2_Plus_TPROJ_FromPlus_L4D3_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_number),
.read_add(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_read_add),
.data_out(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Minus_TPROJ_FromMinus_L4D3_L1L2;
wire PT_L1L2_Minus_TPROJ_FromMinus_L4D3_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_number;
wire [9:0] TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2;
TrackletProjections  TPROJ_FromMinus_L4D3_L1L2(
.data_in(PT_L1L2_Minus_TPROJ_FromMinus_L4D3_L1L2),
.enable(PT_L1L2_Minus_TPROJ_FromMinus_L4D3_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_number),
.read_add(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_read_add),
.data_out(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L4D3(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3_wr_en),
.number_out(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D3;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D3_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L4D3(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D3),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D3_wr_en),
.number_out(TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D3;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D3_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L4D3(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D3),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D3_wr_en),
.number_out(TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Plus_TPROJ_FromPlus_L4D4_L1L2;
wire PT_L1L2_Plus_TPROJ_FromPlus_L4D4_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2;
TrackletProjections  TPROJ_FromPlus_L4D4_L1L2(
.data_in(PT_L1L2_Plus_TPROJ_FromPlus_L4D4_L1L2),
.enable(PT_L1L2_Plus_TPROJ_FromPlus_L4D4_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_number),
.read_add(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Minus_TPROJ_FromMinus_L4D4_L1L2;
wire PT_L1L2_Minus_TPROJ_FromMinus_L4D4_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2;
TrackletProjections  TPROJ_FromMinus_L4D4_L1L2(
.data_in(PT_L1L2_Minus_TPROJ_FromMinus_L4D4_L1L2),
.enable(PT_L1L2_Minus_TPROJ_FromMinus_L4D4_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_number),
.read_add(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L4D4(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4_wr_en),
.number_out(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L4D4(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4_wr_en),
.number_out(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D4;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D4_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L4D4(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D4),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D4_wr_en),
.number_out(TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Plus_TPROJ_FromPlus_L5D3_L1L2;
wire PT_L1L2_Plus_TPROJ_FromPlus_L5D3_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_number;
wire [9:0] TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2;
TrackletProjections  TPROJ_FromPlus_L5D3_L1L2(
.data_in(PT_L1L2_Plus_TPROJ_FromPlus_L5D3_L1L2),
.enable(PT_L1L2_Plus_TPROJ_FromPlus_L5D3_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_number),
.read_add(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_read_add),
.data_out(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Minus_TPROJ_FromMinus_L5D3_L1L2;
wire PT_L1L2_Minus_TPROJ_FromMinus_L5D3_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_number;
wire [9:0] TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2;
TrackletProjections  TPROJ_FromMinus_L5D3_L1L2(
.data_in(PT_L1L2_Minus_TPROJ_FromMinus_L5D3_L1L2),
.enable(PT_L1L2_Minus_TPROJ_FromMinus_L5D3_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_number),
.read_add(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_read_add),
.data_out(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L5D3(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3_wr_en),
.number_out(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D3;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D3_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L5D3(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D3),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D3_wr_en),
.number_out(TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D3;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D3_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L5D3(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D3),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D3_wr_en),
.number_out(TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Plus_TPROJ_FromPlus_L5D4_L1L2;
wire PT_L1L2_Plus_TPROJ_FromPlus_L5D4_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_number;
wire [9:0] TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2;
TrackletProjections  TPROJ_FromPlus_L5D4_L1L2(
.data_in(PT_L1L2_Plus_TPROJ_FromPlus_L5D4_L1L2),
.enable(PT_L1L2_Plus_TPROJ_FromPlus_L5D4_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_number),
.read_add(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_read_add),
.data_out(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Minus_TPROJ_FromMinus_L5D4_L1L2;
wire PT_L1L2_Minus_TPROJ_FromMinus_L5D4_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_number;
wire [9:0] TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2;
TrackletProjections  TPROJ_FromMinus_L5D4_L1L2(
.data_in(PT_L1L2_Minus_TPROJ_FromMinus_L5D4_L1L2),
.enable(PT_L1L2_Minus_TPROJ_FromMinus_L5D4_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_number),
.read_add(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_read_add),
.data_out(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L5D4(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4_wr_en),
.number_out(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D4;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D4_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L5D4(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D4),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D4_wr_en),
.number_out(TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D4;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D4_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L5D4(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D4),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D4_wr_en),
.number_out(TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Plus_TPROJ_FromPlus_L6D3_L1L2;
wire PT_L1L2_Plus_TPROJ_FromPlus_L6D3_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_number;
wire [9:0] TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2;
TrackletProjections  TPROJ_FromPlus_L6D3_L1L2(
.data_in(PT_L1L2_Plus_TPROJ_FromPlus_L6D3_L1L2),
.enable(PT_L1L2_Plus_TPROJ_FromPlus_L6D3_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_number),
.read_add(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_read_add),
.data_out(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Minus_TPROJ_FromMinus_L6D3_L1L2;
wire PT_L1L2_Minus_TPROJ_FromMinus_L6D3_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_number;
wire [9:0] TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2;
TrackletProjections  TPROJ_FromMinus_L6D3_L1L2(
.data_in(PT_L1L2_Minus_TPROJ_FromMinus_L6D3_L1L2),
.enable(PT_L1L2_Minus_TPROJ_FromMinus_L6D3_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_number),
.read_add(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_read_add),
.data_out(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L6D3(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3_wr_en),
.number_out(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D3;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D3_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L6D3(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D3),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D3_wr_en),
.number_out(TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D3;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D3_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L6D3(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D3),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D3_wr_en),
.number_out(TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Plus_TPROJ_FromPlus_L6D4_L1L2;
wire PT_L1L2_Plus_TPROJ_FromPlus_L6D4_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_number;
wire [9:0] TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2;
TrackletProjections  TPROJ_FromPlus_L6D4_L1L2(
.data_in(PT_L1L2_Plus_TPROJ_FromPlus_L6D4_L1L2),
.enable(PT_L1L2_Plus_TPROJ_FromPlus_L6D4_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_number),
.read_add(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_read_add),
.data_out(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L1L2_Minus_TPROJ_FromMinus_L6D4_L1L2;
wire PT_L1L2_Minus_TPROJ_FromMinus_L6D4_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_number;
wire [9:0] TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2;
TrackletProjections  TPROJ_FromMinus_L6D4_L1L2(
.data_in(PT_L1L2_Minus_TPROJ_FromMinus_L6D4_L1L2),
.enable(PT_L1L2_Minus_TPROJ_FromMinus_L6D4_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_number),
.read_add(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_read_add),
.data_out(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L6D4(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4_wr_en),
.number_out(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D4;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D4_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L6D4(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D4),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D4_wr_en),
.number_out(TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D4;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D4_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L6D4(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D4),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D4_wr_en),
.number_out(TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Plus_TPROJ_FromPlus_L1D3_L5L6;
wire PT_L5L6_Plus_TPROJ_FromPlus_L1D3_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6;
TrackletProjections  TPROJ_FromPlus_L1D3_L5L6(
.data_in(PT_L5L6_Plus_TPROJ_FromPlus_L1D3_L5L6),
.enable(PT_L5L6_Plus_TPROJ_FromPlus_L1D3_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_number),
.read_add(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Minus_TPROJ_FromMinus_L1D3_L5L6;
wire PT_L5L6_Minus_TPROJ_FromMinus_L1D3_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6;
TrackletProjections  TPROJ_FromMinus_L1D3_L5L6(
.data_in(PT_L5L6_Minus_TPROJ_FromMinus_L1D3_L5L6),
.enable(PT_L5L6_Minus_TPROJ_FromMinus_L1D3_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_number),
.read_add(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L1D3(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3_wr_en),
.number_out(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L1D3(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3_wr_en),
.number_out(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L1D3(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3_wr_en),
.number_out(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Plus_TPROJ_FromPlus_L1D4_L5L6;
wire PT_L5L6_Plus_TPROJ_FromPlus_L1D4_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_number;
wire [9:0] TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6;
TrackletProjections  TPROJ_FromPlus_L1D4_L5L6(
.data_in(PT_L5L6_Plus_TPROJ_FromPlus_L1D4_L5L6),
.enable(PT_L5L6_Plus_TPROJ_FromPlus_L1D4_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_number),
.read_add(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_read_add),
.data_out(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Minus_TPROJ_FromMinus_L1D4_L5L6;
wire PT_L5L6_Minus_TPROJ_FromMinus_L1D4_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_number;
wire [9:0] TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6;
TrackletProjections  TPROJ_FromMinus_L1D4_L5L6(
.data_in(PT_L5L6_Minus_TPROJ_FromMinus_L1D4_L5L6),
.enable(PT_L5L6_Minus_TPROJ_FromMinus_L1D4_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_number),
.read_add(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_read_add),
.data_out(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D4;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D4_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L1D4(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D4),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D4_wr_en),
.number_out(TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D4;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D4_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L1D4(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D4),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D4_wr_en),
.number_out(TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D4;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D4_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L1D4(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D4),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D4_wr_en),
.number_out(TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Plus_TPROJ_FromPlus_L2D3_L5L6;
wire PT_L5L6_Plus_TPROJ_FromPlus_L2D3_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6;
TrackletProjections  TPROJ_FromPlus_L2D3_L5L6(
.data_in(PT_L5L6_Plus_TPROJ_FromPlus_L2D3_L5L6),
.enable(PT_L5L6_Plus_TPROJ_FromPlus_L2D3_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_number),
.read_add(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Minus_TPROJ_FromMinus_L2D3_L5L6;
wire PT_L5L6_Minus_TPROJ_FromMinus_L2D3_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6;
TrackletProjections  TPROJ_FromMinus_L2D3_L5L6(
.data_in(PT_L5L6_Minus_TPROJ_FromMinus_L2D3_L5L6),
.enable(PT_L5L6_Minus_TPROJ_FromMinus_L2D3_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_number),
.read_add(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L2D3(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3_wr_en),
.number_out(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L2D3(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3_wr_en),
.number_out(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L2D3(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3_wr_en),
.number_out(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Plus_TPROJ_FromPlus_L2D4_L5L6;
wire PT_L5L6_Plus_TPROJ_FromPlus_L2D4_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_number;
wire [9:0] TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6;
TrackletProjections  TPROJ_FromPlus_L2D4_L5L6(
.data_in(PT_L5L6_Plus_TPROJ_FromPlus_L2D4_L5L6),
.enable(PT_L5L6_Plus_TPROJ_FromPlus_L2D4_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_number),
.read_add(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_read_add),
.data_out(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Minus_TPROJ_FromMinus_L2D4_L5L6;
wire PT_L5L6_Minus_TPROJ_FromMinus_L2D4_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_number;
wire [9:0] TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6;
TrackletProjections  TPROJ_FromMinus_L2D4_L5L6(
.data_in(PT_L5L6_Minus_TPROJ_FromMinus_L2D4_L5L6),
.enable(PT_L5L6_Minus_TPROJ_FromMinus_L2D4_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_number),
.read_add(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_read_add),
.data_out(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D4;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D4_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L2D4(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D4),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D4_wr_en),
.number_out(TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D4;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D4_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L2D4(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D4),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D4_wr_en),
.number_out(TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D4;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D4_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L2D4(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D4),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D4_wr_en),
.number_out(TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Plus_TPROJ_FromPlus_L3D3_L5L6;
wire PT_L5L6_Plus_TPROJ_FromPlus_L3D3_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6;
TrackletProjections  TPROJ_FromPlus_L3D3_L5L6(
.data_in(PT_L5L6_Plus_TPROJ_FromPlus_L3D3_L5L6),
.enable(PT_L5L6_Plus_TPROJ_FromPlus_L3D3_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_number),
.read_add(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Minus_TPROJ_FromMinus_L3D3_L5L6;
wire PT_L5L6_Minus_TPROJ_FromMinus_L3D3_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6;
TrackletProjections  TPROJ_FromMinus_L3D3_L5L6(
.data_in(PT_L5L6_Minus_TPROJ_FromMinus_L3D3_L5L6),
.enable(PT_L5L6_Minus_TPROJ_FromMinus_L3D3_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_number),
.read_add(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L3D3(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3_wr_en),
.number_out(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L3D3(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3_wr_en),
.number_out(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L3D3(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3_wr_en),
.number_out(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Plus_TPROJ_FromPlus_L3D4_L5L6;
wire PT_L5L6_Plus_TPROJ_FromPlus_L3D4_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_number;
wire [9:0] TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6;
TrackletProjections  TPROJ_FromPlus_L3D4_L5L6(
.data_in(PT_L5L6_Plus_TPROJ_FromPlus_L3D4_L5L6),
.enable(PT_L5L6_Plus_TPROJ_FromPlus_L3D4_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_number),
.read_add(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_read_add),
.data_out(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Minus_TPROJ_FromMinus_L3D4_L5L6;
wire PT_L5L6_Minus_TPROJ_FromMinus_L3D4_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_number;
wire [9:0] TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6;
TrackletProjections  TPROJ_FromMinus_L3D4_L5L6(
.data_in(PT_L5L6_Minus_TPROJ_FromMinus_L3D4_L5L6),
.enable(PT_L5L6_Minus_TPROJ_FromMinus_L3D4_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_number),
.read_add(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_read_add),
.data_out(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D4;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D4_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L3D4(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D4),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D4_wr_en),
.number_out(TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D4;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D4_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L3D4(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D4),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D4_wr_en),
.number_out(TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L3D4(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4_wr_en),
.number_out(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Plus_TPROJ_FromPlus_L4D3_L5L6;
wire PT_L5L6_Plus_TPROJ_FromPlus_L4D3_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6;
TrackletProjections  TPROJ_FromPlus_L4D3_L5L6(
.data_in(PT_L5L6_Plus_TPROJ_FromPlus_L4D3_L5L6),
.enable(PT_L5L6_Plus_TPROJ_FromPlus_L4D3_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_number),
.read_add(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Minus_TPROJ_FromMinus_L4D3_L5L6;
wire PT_L5L6_Minus_TPROJ_FromMinus_L4D3_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6;
TrackletProjections  TPROJ_FromMinus_L4D3_L5L6(
.data_in(PT_L5L6_Minus_TPROJ_FromMinus_L4D3_L5L6),
.enable(PT_L5L6_Minus_TPROJ_FromMinus_L4D3_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_number),
.read_add(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L4D3(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3_wr_en),
.number_out(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L4D3(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3_wr_en),
.number_out(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L4D3(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3_wr_en),
.number_out(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Plus_TPROJ_FromPlus_L4D4_L5L6;
wire PT_L5L6_Plus_TPROJ_FromPlus_L4D4_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_number;
wire [9:0] TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6;
TrackletProjections  TPROJ_FromPlus_L4D4_L5L6(
.data_in(PT_L5L6_Plus_TPROJ_FromPlus_L4D4_L5L6),
.enable(PT_L5L6_Plus_TPROJ_FromPlus_L4D4_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_number),
.read_add(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_read_add),
.data_out(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] PT_L5L6_Minus_TPROJ_FromMinus_L4D4_L5L6;
wire PT_L5L6_Minus_TPROJ_FromMinus_L4D4_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_number;
wire [9:0] TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6;
TrackletProjections  TPROJ_FromMinus_L4D4_L5L6(
.data_in(PT_L5L6_Minus_TPROJ_FromMinus_L4D4_L5L6),
.enable(PT_L5L6_Minus_TPROJ_FromMinus_L4D4_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_number),
.read_add(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_read_add),
.data_out(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6),
.start(start6_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D4;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D4_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L4D4(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D4),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D4_wr_en),
.number_out(TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D4;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D4_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L4D4(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D4),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D4_wr_en),
.number_out(TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L4D4(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4_wr_en),
.number_out(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6),
.start(startproj5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z1;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1;
VMProjections  VMPROJ_L3L4_L1D3PHI1Z1(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z1),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z1_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1_number),
.read_add(VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1),
.start(start7_0),
.done(done6_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z1n7;
wire VMR_L1D3_VMS_L1D3PHI1Z1n7_wr_en;
wire [5:0] VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1_number;
wire [10:0] VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1_read_add;
wire [17:0] VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1;
VMStubs #("Match") VMS_L1D3PHI1Z1n7(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z1n7),
.enable(VMR_L1D3_VMS_L1D3PHI1Z1n7_wr_en),
.number_out(VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1_number),
.read_add(VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1_read_add),
.data_out(VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z2;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2;
VMProjections  VMPROJ_L3L4_L1D3PHI1Z2(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z2),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z2_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2_number),
.read_add(VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z2n7;
wire VMR_L1D3_VMS_L1D3PHI1Z2n7_wr_en;
wire [5:0] VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2_number;
wire [10:0] VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2_read_add;
wire [17:0] VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2;
VMStubs #("Match") VMS_L1D3PHI1Z2n7(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z2n7),
.enable(VMR_L1D3_VMS_L1D3PHI1Z2n7_wr_en),
.number_out(VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2_number),
.read_add(VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2_read_add),
.data_out(VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z1;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1;
VMProjections  VMPROJ_L3L4_L1D3PHI2Z1(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z1),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z1_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1_number),
.read_add(VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z1n7;
wire VMR_L1D3_VMS_L1D3PHI2Z1n7_wr_en;
wire [5:0] VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1_number;
wire [10:0] VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1_read_add;
wire [17:0] VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1;
VMStubs #("Match") VMS_L1D3PHI2Z1n7(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z1n7),
.enable(VMR_L1D3_VMS_L1D3PHI2Z1n7_wr_en),
.number_out(VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1_number),
.read_add(VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1_read_add),
.data_out(VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z2;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2;
VMProjections  VMPROJ_L3L4_L1D3PHI2Z2(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z2),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z2_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2_number),
.read_add(VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z2n7;
wire VMR_L1D3_VMS_L1D3PHI2Z2n7_wr_en;
wire [5:0] VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2_number;
wire [10:0] VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2_read_add;
wire [17:0] VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2;
VMStubs #("Match") VMS_L1D3PHI2Z2n7(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z2n7),
.enable(VMR_L1D3_VMS_L1D3PHI2Z2n7_wr_en),
.number_out(VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2_number),
.read_add(VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2_read_add),
.data_out(VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z1;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1;
VMProjections  VMPROJ_L3L4_L1D3PHI3Z1(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z1),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z1_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1_number),
.read_add(VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z1n7;
wire VMR_L1D3_VMS_L1D3PHI3Z1n7_wr_en;
wire [5:0] VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1_number;
wire [10:0] VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1_read_add;
wire [17:0] VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1;
VMStubs #("Match") VMS_L1D3PHI3Z1n7(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z1n7),
.enable(VMR_L1D3_VMS_L1D3PHI3Z1n7_wr_en),
.number_out(VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1_number),
.read_add(VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1_read_add),
.data_out(VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z2;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2;
VMProjections  VMPROJ_L3L4_L1D3PHI3Z2(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z2),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z2_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2_number),
.read_add(VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z2n7;
wire VMR_L1D3_VMS_L1D3PHI3Z2n7_wr_en;
wire [5:0] VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2_number;
wire [10:0] VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2_read_add;
wire [17:0] VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2;
VMStubs #("Match") VMS_L1D3PHI3Z2n7(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z2n7),
.enable(VMR_L1D3_VMS_L1D3PHI3Z2n7_wr_en),
.number_out(VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2_number),
.read_add(VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2_read_add),
.data_out(VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z1;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1;
VMProjections  VMPROJ_L3L4_L1D4PHI1Z1(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z1),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z1_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1_number),
.read_add(VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI1Z1n3;
wire VMR_L1D4_VMS_L1D4PHI1Z1n3_wr_en;
wire [5:0] VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1_number;
wire [10:0] VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1_read_add;
wire [17:0] VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1;
VMStubs #("Match") VMS_L1D4PHI1Z1n3(
.data_in(VMR_L1D4_VMS_L1D4PHI1Z1n3),
.enable(VMR_L1D4_VMS_L1D4PHI1Z1n3_wr_en),
.number_out(VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1_number),
.read_add(VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1_read_add),
.data_out(VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z2;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2;
VMProjections  VMPROJ_L3L4_L1D4PHI1Z2(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z2),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z2_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2_number),
.read_add(VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI1Z2n1;
wire VMR_L1D4_VMS_L1D4PHI1Z2n1_wr_en;
wire [5:0] VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2_number;
wire [10:0] VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2_read_add;
wire [17:0] VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2;
VMStubs #("Match") VMS_L1D4PHI1Z2n1(
.data_in(VMR_L1D4_VMS_L1D4PHI1Z2n1),
.enable(VMR_L1D4_VMS_L1D4PHI1Z2n1_wr_en),
.number_out(VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2_number),
.read_add(VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2_read_add),
.data_out(VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z1;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1;
VMProjections  VMPROJ_L3L4_L1D4PHI2Z1(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z1),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z1_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1_number),
.read_add(VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI2Z1n3;
wire VMR_L1D4_VMS_L1D4PHI2Z1n3_wr_en;
wire [5:0] VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1_number;
wire [10:0] VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1_read_add;
wire [17:0] VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1;
VMStubs #("Match") VMS_L1D4PHI2Z1n3(
.data_in(VMR_L1D4_VMS_L1D4PHI2Z1n3),
.enable(VMR_L1D4_VMS_L1D4PHI2Z1n3_wr_en),
.number_out(VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1_number),
.read_add(VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1_read_add),
.data_out(VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z2;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2;
VMProjections  VMPROJ_L3L4_L1D4PHI2Z2(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z2),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z2_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2_number),
.read_add(VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI2Z2n1;
wire VMR_L1D4_VMS_L1D4PHI2Z2n1_wr_en;
wire [5:0] VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2_number;
wire [10:0] VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2_read_add;
wire [17:0] VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2;
VMStubs #("Match") VMS_L1D4PHI2Z2n1(
.data_in(VMR_L1D4_VMS_L1D4PHI2Z2n1),
.enable(VMR_L1D4_VMS_L1D4PHI2Z2n1_wr_en),
.number_out(VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2_number),
.read_add(VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2_read_add),
.data_out(VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z1;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1;
VMProjections  VMPROJ_L3L4_L1D4PHI3Z1(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z1),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z1_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1_number),
.read_add(VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI3Z1n3;
wire VMR_L1D4_VMS_L1D4PHI3Z1n3_wr_en;
wire [5:0] VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1_number;
wire [10:0] VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1_read_add;
wire [17:0] VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1;
VMStubs #("Match") VMS_L1D4PHI3Z1n3(
.data_in(VMR_L1D4_VMS_L1D4PHI3Z1n3),
.enable(VMR_L1D4_VMS_L1D4PHI3Z1n3_wr_en),
.number_out(VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1_number),
.read_add(VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1_read_add),
.data_out(VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z2;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2;
VMProjections  VMPROJ_L3L4_L1D4PHI3Z2(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z2),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z2_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2_number),
.read_add(VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI3Z2n1;
wire VMR_L1D4_VMS_L1D4PHI3Z2n1_wr_en;
wire [5:0] VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2_number;
wire [10:0] VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2_read_add;
wire [17:0] VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2;
VMStubs #("Match") VMS_L1D4PHI3Z2n1(
.data_in(VMR_L1D4_VMS_L1D4PHI3Z2n1),
.enable(VMR_L1D4_VMS_L1D4PHI3Z2n1_wr_en),
.number_out(VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2_number),
.read_add(VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2_read_add),
.data_out(VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z1;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1;
VMProjections  VMPROJ_L3L4_L2D3PHI1Z1(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z1),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z1_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1_number),
.read_add(VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI1Z1n2;
wire VMR_L2D3_VMS_L2D3PHI1Z1n2_wr_en;
wire [5:0] VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1_number;
wire [10:0] VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1_read_add;
wire [17:0] VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1;
VMStubs #("Match") VMS_L2D3PHI1Z1n2(
.data_in(VMR_L2D3_VMS_L2D3PHI1Z1n2),
.enable(VMR_L2D3_VMS_L2D3PHI1Z1n2_wr_en),
.number_out(VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1_number),
.read_add(VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1_read_add),
.data_out(VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z2;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2;
VMProjections  VMPROJ_L3L4_L2D3PHI1Z2(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z2),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z2_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2_number),
.read_add(VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI1Z2n3;
wire VMR_L2D3_VMS_L2D3PHI1Z2n3_wr_en;
wire [5:0] VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2_number;
wire [10:0] VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2_read_add;
wire [17:0] VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2;
VMStubs #("Match") VMS_L2D3PHI1Z2n3(
.data_in(VMR_L2D3_VMS_L2D3PHI1Z2n3),
.enable(VMR_L2D3_VMS_L2D3PHI1Z2n3_wr_en),
.number_out(VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2_number),
.read_add(VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2_read_add),
.data_out(VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z1;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1;
VMProjections  VMPROJ_L3L4_L2D3PHI2Z1(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z1),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z1_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1_number),
.read_add(VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z1n3;
wire VMR_L2D3_VMS_L2D3PHI2Z1n3_wr_en;
wire [5:0] VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1_number;
wire [10:0] VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1_read_add;
wire [17:0] VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1;
VMStubs #("Match") VMS_L2D3PHI2Z1n3(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z1n3),
.enable(VMR_L2D3_VMS_L2D3PHI2Z1n3_wr_en),
.number_out(VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1_number),
.read_add(VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1_read_add),
.data_out(VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z2;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2;
VMProjections  VMPROJ_L3L4_L2D3PHI2Z2(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z2),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z2_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2_number),
.read_add(VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z2n5;
wire VMR_L2D3_VMS_L2D3PHI2Z2n5_wr_en;
wire [5:0] VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2_number;
wire [10:0] VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2;
VMStubs #("Match") VMS_L2D3PHI2Z2n5(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z2n5),
.enable(VMR_L2D3_VMS_L2D3PHI2Z2n5_wr_en),
.number_out(VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2_number),
.read_add(VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2_read_add),
.data_out(VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z1;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1;
VMProjections  VMPROJ_L3L4_L2D3PHI3Z1(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z1),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z1_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1_number),
.read_add(VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z1n3;
wire VMR_L2D3_VMS_L2D3PHI3Z1n3_wr_en;
wire [5:0] VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1_number;
wire [10:0] VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1_read_add;
wire [17:0] VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1;
VMStubs #("Match") VMS_L2D3PHI3Z1n3(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z1n3),
.enable(VMR_L2D3_VMS_L2D3PHI3Z1n3_wr_en),
.number_out(VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1_number),
.read_add(VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1_read_add),
.data_out(VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z2;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2;
VMProjections  VMPROJ_L3L4_L2D3PHI3Z2(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z2),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z2_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2_number),
.read_add(VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z2n5;
wire VMR_L2D3_VMS_L2D3PHI3Z2n5_wr_en;
wire [5:0] VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2_number;
wire [10:0] VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2;
VMStubs #("Match") VMS_L2D3PHI3Z2n5(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z2n5),
.enable(VMR_L2D3_VMS_L2D3PHI3Z2n5_wr_en),
.number_out(VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2_number),
.read_add(VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2_read_add),
.data_out(VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z1;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1_read_add;
wire [12:0] VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1;
VMProjections  VMPROJ_L3L4_L2D3PHI4Z1(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z1),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z1_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1_number),
.read_add(VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI4Z1n2;
wire VMR_L2D3_VMS_L2D3PHI4Z1n2_wr_en;
wire [5:0] VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1_number;
wire [10:0] VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1_read_add;
wire [17:0] VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1;
VMStubs #("Match") VMS_L2D3PHI4Z1n2(
.data_in(VMR_L2D3_VMS_L2D3PHI4Z1n2),
.enable(VMR_L2D3_VMS_L2D3PHI4Z1n2_wr_en),
.number_out(VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1_number),
.read_add(VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1_read_add),
.data_out(VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z2;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2_read_add;
wire [12:0] VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2;
VMProjections  VMPROJ_L3L4_L2D3PHI4Z2(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z2),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z2_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2_number),
.read_add(VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI4Z2n3;
wire VMR_L2D3_VMS_L2D3PHI4Z2n3_wr_en;
wire [5:0] VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2_number;
wire [10:0] VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2_read_add;
wire [17:0] VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2;
VMStubs #("Match") VMS_L2D3PHI4Z2n3(
.data_in(VMR_L2D3_VMS_L2D3PHI4Z2n3),
.enable(VMR_L2D3_VMS_L2D3PHI4Z2n3_wr_en),
.number_out(VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2_number),
.read_add(VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2_read_add),
.data_out(VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z1;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1;
VMProjections  VMPROJ_L3L4_L2D4PHI1Z1(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z1),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z1_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1_number),
.read_add(VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI1Z1n3;
wire VMR_L2D4_VMS_L2D4PHI1Z1n3_wr_en;
wire [5:0] VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1_number;
wire [10:0] VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1_read_add;
wire [17:0] VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1;
VMStubs #("Match") VMS_L2D4PHI1Z1n3(
.data_in(VMR_L2D4_VMS_L2D4PHI1Z1n3),
.enable(VMR_L2D4_VMS_L2D4PHI1Z1n3_wr_en),
.number_out(VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1_number),
.read_add(VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1_read_add),
.data_out(VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z2;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2;
VMProjections  VMPROJ_L3L4_L2D4PHI1Z2(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z2),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z2_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2_number),
.read_add(VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI1Z2n3;
wire VMR_L2D4_VMS_L2D4PHI1Z2n3_wr_en;
wire [5:0] VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2_number;
wire [10:0] VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2_read_add;
wire [17:0] VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2;
VMStubs #("Match") VMS_L2D4PHI1Z2n3(
.data_in(VMR_L2D4_VMS_L2D4PHI1Z2n3),
.enable(VMR_L2D4_VMS_L2D4PHI1Z2n3_wr_en),
.number_out(VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2_number),
.read_add(VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2_read_add),
.data_out(VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z1;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1;
VMProjections  VMPROJ_L3L4_L2D4PHI2Z1(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z1),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z1_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1_number),
.read_add(VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z1n5;
wire VMR_L2D4_VMS_L2D4PHI2Z1n5_wr_en;
wire [5:0] VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1_number;
wire [10:0] VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1;
VMStubs #("Match") VMS_L2D4PHI2Z1n5(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z1n5),
.enable(VMR_L2D4_VMS_L2D4PHI2Z1n5_wr_en),
.number_out(VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1_number),
.read_add(VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1_read_add),
.data_out(VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z2;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2;
VMProjections  VMPROJ_L3L4_L2D4PHI2Z2(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z2),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z2_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2_number),
.read_add(VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z2n5;
wire VMR_L2D4_VMS_L2D4PHI2Z2n5_wr_en;
wire [5:0] VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2_number;
wire [10:0] VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2;
VMStubs #("Match") VMS_L2D4PHI2Z2n5(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z2n5),
.enable(VMR_L2D4_VMS_L2D4PHI2Z2n5_wr_en),
.number_out(VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2_number),
.read_add(VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2_read_add),
.data_out(VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z1;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1;
VMProjections  VMPROJ_L3L4_L2D4PHI3Z1(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z1),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z1_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1_number),
.read_add(VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z1n5;
wire VMR_L2D4_VMS_L2D4PHI3Z1n5_wr_en;
wire [5:0] VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1_number;
wire [10:0] VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1;
VMStubs #("Match") VMS_L2D4PHI3Z1n5(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z1n5),
.enable(VMR_L2D4_VMS_L2D4PHI3Z1n5_wr_en),
.number_out(VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1_number),
.read_add(VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1_read_add),
.data_out(VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z2;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2;
VMProjections  VMPROJ_L3L4_L2D4PHI3Z2(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z2),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z2_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2_number),
.read_add(VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z2n5;
wire VMR_L2D4_VMS_L2D4PHI3Z2n5_wr_en;
wire [5:0] VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2_number;
wire [10:0] VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2;
VMStubs #("Match") VMS_L2D4PHI3Z2n5(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z2n5),
.enable(VMR_L2D4_VMS_L2D4PHI3Z2n5_wr_en),
.number_out(VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2_number),
.read_add(VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2_read_add),
.data_out(VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z1;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1_read_add;
wire [12:0] VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1;
VMProjections  VMPROJ_L3L4_L2D4PHI4Z1(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z1),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z1_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1_number),
.read_add(VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI4Z1n3;
wire VMR_L2D4_VMS_L2D4PHI4Z1n3_wr_en;
wire [5:0] VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1_number;
wire [10:0] VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1_read_add;
wire [17:0] VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1;
VMStubs #("Match") VMS_L2D4PHI4Z1n3(
.data_in(VMR_L2D4_VMS_L2D4PHI4Z1n3),
.enable(VMR_L2D4_VMS_L2D4PHI4Z1n3_wr_en),
.number_out(VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1_number),
.read_add(VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1_read_add),
.data_out(VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z2;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2_read_add;
wire [12:0] VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2;
VMProjections  VMPROJ_L3L4_L2D4PHI4Z2(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z2),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z2_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2_number),
.read_add(VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI4Z2n3;
wire VMR_L2D4_VMS_L2D4PHI4Z2n3_wr_en;
wire [5:0] VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2_number;
wire [10:0] VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2_read_add;
wire [17:0] VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2;
VMStubs #("Match") VMS_L2D4PHI4Z2n3(
.data_in(VMR_L2D4_VMS_L2D4PHI4Z2n3),
.enable(VMR_L2D4_VMS_L2D4PHI4Z2n3_wr_en),
.number_out(VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2_number),
.read_add(VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2_read_add),
.data_out(VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z1;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1;
VMProjections  VMPROJ_L3L4_L5D3PHI1Z1(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z1),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z1_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1_number),
.read_add(VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z1n5;
wire VMR_L5D3_VMS_L5D3PHI1Z1n5_wr_en;
wire [5:0] VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1_number;
wire [10:0] VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1_read_add;
wire [17:0] VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1;
VMStubs #("Match") VMS_L5D3PHI1Z1n5(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z1n5),
.enable(VMR_L5D3_VMS_L5D3PHI1Z1n5_wr_en),
.number_out(VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1_number),
.read_add(VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1_read_add),
.data_out(VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z2;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2;
VMProjections  VMPROJ_L3L4_L5D3PHI1Z2(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z2),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z2_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2_number),
.read_add(VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z2n5;
wire VMR_L5D3_VMS_L5D3PHI1Z2n5_wr_en;
wire [5:0] VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2_number;
wire [10:0] VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2_read_add;
wire [17:0] VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2;
VMStubs #("Match") VMS_L5D3PHI1Z2n5(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z2n5),
.enable(VMR_L5D3_VMS_L5D3PHI1Z2n5_wr_en),
.number_out(VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2_number),
.read_add(VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2_read_add),
.data_out(VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z1;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1;
VMProjections  VMPROJ_L3L4_L5D3PHI2Z1(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z1),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z1_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1_number),
.read_add(VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z1n5;
wire VMR_L5D3_VMS_L5D3PHI2Z1n5_wr_en;
wire [5:0] VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1_number;
wire [10:0] VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1_read_add;
wire [17:0] VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1;
VMStubs #("Match") VMS_L5D3PHI2Z1n5(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z1n5),
.enable(VMR_L5D3_VMS_L5D3PHI2Z1n5_wr_en),
.number_out(VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1_number),
.read_add(VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1_read_add),
.data_out(VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z2;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2;
VMProjections  VMPROJ_L3L4_L5D3PHI2Z2(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z2),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z2_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2_number),
.read_add(VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z2n5;
wire VMR_L5D3_VMS_L5D3PHI2Z2n5_wr_en;
wire [5:0] VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2_number;
wire [10:0] VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2_read_add;
wire [17:0] VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2;
VMStubs #("Match") VMS_L5D3PHI2Z2n5(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z2n5),
.enable(VMR_L5D3_VMS_L5D3PHI2Z2n5_wr_en),
.number_out(VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2_number),
.read_add(VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2_read_add),
.data_out(VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z1;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1;
VMProjections  VMPROJ_L3L4_L5D3PHI3Z1(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z1),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z1_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1_number),
.read_add(VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z1n5;
wire VMR_L5D3_VMS_L5D3PHI3Z1n5_wr_en;
wire [5:0] VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1_number;
wire [10:0] VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1_read_add;
wire [17:0] VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1;
VMStubs #("Match") VMS_L5D3PHI3Z1n5(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z1n5),
.enable(VMR_L5D3_VMS_L5D3PHI3Z1n5_wr_en),
.number_out(VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1_number),
.read_add(VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1_read_add),
.data_out(VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z2;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2;
VMProjections  VMPROJ_L3L4_L5D3PHI3Z2(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z2),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z2_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2_number),
.read_add(VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z2n5;
wire VMR_L5D3_VMS_L5D3PHI3Z2n5_wr_en;
wire [5:0] VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2_number;
wire [10:0] VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2_read_add;
wire [17:0] VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2;
VMStubs #("Match") VMS_L5D3PHI3Z2n5(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z2n5),
.enable(VMR_L5D3_VMS_L5D3PHI3Z2n5_wr_en),
.number_out(VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2_number),
.read_add(VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2_read_add),
.data_out(VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z1;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1;
VMProjections  VMPROJ_L3L4_L5D4PHI1Z1(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z1),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z1_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1_number),
.read_add(VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z1n5;
wire VMR_L5D4_VMS_L5D4PHI1Z1n5_wr_en;
wire [5:0] VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1_number;
wire [10:0] VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1_read_add;
wire [17:0] VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1;
VMStubs #("Match") VMS_L5D4PHI1Z1n5(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z1n5),
.enable(VMR_L5D4_VMS_L5D4PHI1Z1n5_wr_en),
.number_out(VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1_number),
.read_add(VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1_read_add),
.data_out(VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z2;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2;
VMProjections  VMPROJ_L3L4_L5D4PHI1Z2(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z2),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z2_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2_number),
.read_add(VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z2n3;
wire VMR_L5D4_VMS_L5D4PHI1Z2n3_wr_en;
wire [5:0] VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2_number;
wire [10:0] VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2_read_add;
wire [17:0] VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2;
VMStubs #("Match") VMS_L5D4PHI1Z2n3(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z2n3),
.enable(VMR_L5D4_VMS_L5D4PHI1Z2n3_wr_en),
.number_out(VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2_number),
.read_add(VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2_read_add),
.data_out(VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z1;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1;
VMProjections  VMPROJ_L3L4_L5D4PHI2Z1(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z1),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z1_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1_number),
.read_add(VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z1n5;
wire VMR_L5D4_VMS_L5D4PHI2Z1n5_wr_en;
wire [5:0] VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1_number;
wire [10:0] VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1_read_add;
wire [17:0] VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1;
VMStubs #("Match") VMS_L5D4PHI2Z1n5(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z1n5),
.enable(VMR_L5D4_VMS_L5D4PHI2Z1n5_wr_en),
.number_out(VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1_number),
.read_add(VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1_read_add),
.data_out(VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z2;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2;
VMProjections  VMPROJ_L3L4_L5D4PHI2Z2(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z2),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z2_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2_number),
.read_add(VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z2n3;
wire VMR_L5D4_VMS_L5D4PHI2Z2n3_wr_en;
wire [5:0] VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2_number;
wire [10:0] VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2_read_add;
wire [17:0] VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2;
VMStubs #("Match") VMS_L5D4PHI2Z2n3(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z2n3),
.enable(VMR_L5D4_VMS_L5D4PHI2Z2n3_wr_en),
.number_out(VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2_number),
.read_add(VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2_read_add),
.data_out(VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z1;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1;
VMProjections  VMPROJ_L3L4_L5D4PHI3Z1(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z1),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z1_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1_number),
.read_add(VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z1n5;
wire VMR_L5D4_VMS_L5D4PHI3Z1n5_wr_en;
wire [5:0] VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1_number;
wire [10:0] VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1_read_add;
wire [17:0] VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1;
VMStubs #("Match") VMS_L5D4PHI3Z1n5(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z1n5),
.enable(VMR_L5D4_VMS_L5D4PHI3Z1n5_wr_en),
.number_out(VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1_number),
.read_add(VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1_read_add),
.data_out(VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z2;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2;
VMProjections  VMPROJ_L3L4_L5D4PHI3Z2(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z2),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z2_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2_number),
.read_add(VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z2n3;
wire VMR_L5D4_VMS_L5D4PHI3Z2n3_wr_en;
wire [5:0] VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2_number;
wire [10:0] VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2_read_add;
wire [17:0] VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2;
VMStubs #("Match") VMS_L5D4PHI3Z2n3(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z2n3),
.enable(VMR_L5D4_VMS_L5D4PHI3Z2n3_wr_en),
.number_out(VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2_number),
.read_add(VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2_read_add),
.data_out(VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z1;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1;
VMProjections  VMPROJ_L3L4_L6D3PHI1Z1(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z1),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z1_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1_number),
.read_add(VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI1Z1n2;
wire VMR_L6D3_VMS_L6D3PHI1Z1n2_wr_en;
wire [5:0] VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1_number;
wire [10:0] VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1_read_add;
wire [17:0] VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1;
VMStubs #("Match") VMS_L6D3PHI1Z1n2(
.data_in(VMR_L6D3_VMS_L6D3PHI1Z1n2),
.enable(VMR_L6D3_VMS_L6D3PHI1Z1n2_wr_en),
.number_out(VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1_number),
.read_add(VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1_read_add),
.data_out(VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z2;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2;
VMProjections  VMPROJ_L3L4_L6D3PHI1Z2(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z2),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z2_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2_number),
.read_add(VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI1Z2n3;
wire VMR_L6D3_VMS_L6D3PHI1Z2n3_wr_en;
wire [5:0] VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2_number;
wire [10:0] VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2_read_add;
wire [17:0] VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2;
VMStubs #("Match") VMS_L6D3PHI1Z2n3(
.data_in(VMR_L6D3_VMS_L6D3PHI1Z2n3),
.enable(VMR_L6D3_VMS_L6D3PHI1Z2n3_wr_en),
.number_out(VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2_number),
.read_add(VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2_read_add),
.data_out(VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z1;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1;
VMProjections  VMPROJ_L3L4_L6D3PHI2Z1(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z1),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z1_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1_number),
.read_add(VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z1n3;
wire VMR_L6D3_VMS_L6D3PHI2Z1n3_wr_en;
wire [5:0] VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1_number;
wire [10:0] VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1_read_add;
wire [17:0] VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1;
VMStubs #("Match") VMS_L6D3PHI2Z1n3(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z1n3),
.enable(VMR_L6D3_VMS_L6D3PHI2Z1n3_wr_en),
.number_out(VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1_number),
.read_add(VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1_read_add),
.data_out(VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z2;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2;
VMProjections  VMPROJ_L3L4_L6D3PHI2Z2(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z2),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z2_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2_number),
.read_add(VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z2n5;
wire VMR_L6D3_VMS_L6D3PHI2Z2n5_wr_en;
wire [5:0] VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2_number;
wire [10:0] VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2;
VMStubs #("Match") VMS_L6D3PHI2Z2n5(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z2n5),
.enable(VMR_L6D3_VMS_L6D3PHI2Z2n5_wr_en),
.number_out(VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2_number),
.read_add(VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2_read_add),
.data_out(VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z1;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1;
VMProjections  VMPROJ_L3L4_L6D3PHI3Z1(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z1),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z1_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1_number),
.read_add(VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z1n3;
wire VMR_L6D3_VMS_L6D3PHI3Z1n3_wr_en;
wire [5:0] VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1_number;
wire [10:0] VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1_read_add;
wire [17:0] VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1;
VMStubs #("Match") VMS_L6D3PHI3Z1n3(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z1n3),
.enable(VMR_L6D3_VMS_L6D3PHI3Z1n3_wr_en),
.number_out(VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1_number),
.read_add(VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1_read_add),
.data_out(VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z2;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2;
VMProjections  VMPROJ_L3L4_L6D3PHI3Z2(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z2),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z2_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2_number),
.read_add(VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z2n5;
wire VMR_L6D3_VMS_L6D3PHI3Z2n5_wr_en;
wire [5:0] VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2_number;
wire [10:0] VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2;
VMStubs #("Match") VMS_L6D3PHI3Z2n5(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z2n5),
.enable(VMR_L6D3_VMS_L6D3PHI3Z2n5_wr_en),
.number_out(VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2_number),
.read_add(VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2_read_add),
.data_out(VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z1;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1_read_add;
wire [12:0] VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1;
VMProjections  VMPROJ_L3L4_L6D3PHI4Z1(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z1),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z1_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1_number),
.read_add(VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI4Z1n2;
wire VMR_L6D3_VMS_L6D3PHI4Z1n2_wr_en;
wire [5:0] VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1_number;
wire [10:0] VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1_read_add;
wire [17:0] VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1;
VMStubs #("Match") VMS_L6D3PHI4Z1n2(
.data_in(VMR_L6D3_VMS_L6D3PHI4Z1n2),
.enable(VMR_L6D3_VMS_L6D3PHI4Z1n2_wr_en),
.number_out(VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1_number),
.read_add(VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1_read_add),
.data_out(VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z2;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2_read_add;
wire [12:0] VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2;
VMProjections  VMPROJ_L3L4_L6D3PHI4Z2(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z2),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z2_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2_number),
.read_add(VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI4Z2n3;
wire VMR_L6D3_VMS_L6D3PHI4Z2n3_wr_en;
wire [5:0] VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2_number;
wire [10:0] VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2_read_add;
wire [17:0] VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2;
VMStubs #("Match") VMS_L6D3PHI4Z2n3(
.data_in(VMR_L6D3_VMS_L6D3PHI4Z2n3),
.enable(VMR_L6D3_VMS_L6D3PHI4Z2n3_wr_en),
.number_out(VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2_number),
.read_add(VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2_read_add),
.data_out(VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z1;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1;
VMProjections  VMPROJ_L3L4_L6D4PHI1Z1(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z1),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z1_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1_number),
.read_add(VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI1Z1n3;
wire VMR_L6D4_VMS_L6D4PHI1Z1n3_wr_en;
wire [5:0] VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1_number;
wire [10:0] VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1_read_add;
wire [17:0] VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1;
VMStubs #("Match") VMS_L6D4PHI1Z1n3(
.data_in(VMR_L6D4_VMS_L6D4PHI1Z1n3),
.enable(VMR_L6D4_VMS_L6D4PHI1Z1n3_wr_en),
.number_out(VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1_number),
.read_add(VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1_read_add),
.data_out(VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z2;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2;
VMProjections  VMPROJ_L3L4_L6D4PHI1Z2(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z2),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z2_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2_number),
.read_add(VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI1Z2n3;
wire VMR_L6D4_VMS_L6D4PHI1Z2n3_wr_en;
wire [5:0] VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2_number;
wire [10:0] VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2_read_add;
wire [17:0] VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2;
VMStubs #("Match") VMS_L6D4PHI1Z2n3(
.data_in(VMR_L6D4_VMS_L6D4PHI1Z2n3),
.enable(VMR_L6D4_VMS_L6D4PHI1Z2n3_wr_en),
.number_out(VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2_number),
.read_add(VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2_read_add),
.data_out(VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z1;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1;
VMProjections  VMPROJ_L3L4_L6D4PHI2Z1(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z1),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z1_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1_number),
.read_add(VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z1n5;
wire VMR_L6D4_VMS_L6D4PHI2Z1n5_wr_en;
wire [5:0] VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1_number;
wire [10:0] VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1;
VMStubs #("Match") VMS_L6D4PHI2Z1n5(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z1n5),
.enable(VMR_L6D4_VMS_L6D4PHI2Z1n5_wr_en),
.number_out(VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1_number),
.read_add(VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1_read_add),
.data_out(VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z2;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2;
VMProjections  VMPROJ_L3L4_L6D4PHI2Z2(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z2),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z2_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2_number),
.read_add(VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z2n5;
wire VMR_L6D4_VMS_L6D4PHI2Z2n5_wr_en;
wire [5:0] VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2_number;
wire [10:0] VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2;
VMStubs #("Match") VMS_L6D4PHI2Z2n5(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z2n5),
.enable(VMR_L6D4_VMS_L6D4PHI2Z2n5_wr_en),
.number_out(VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2_number),
.read_add(VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2_read_add),
.data_out(VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z1;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1;
VMProjections  VMPROJ_L3L4_L6D4PHI3Z1(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z1),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z1_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1_number),
.read_add(VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z1n5;
wire VMR_L6D4_VMS_L6D4PHI3Z1n5_wr_en;
wire [5:0] VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1_number;
wire [10:0] VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1;
VMStubs #("Match") VMS_L6D4PHI3Z1n5(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z1n5),
.enable(VMR_L6D4_VMS_L6D4PHI3Z1n5_wr_en),
.number_out(VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1_number),
.read_add(VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1_read_add),
.data_out(VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z2;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2;
VMProjections  VMPROJ_L3L4_L6D4PHI3Z2(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z2),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z2_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2_number),
.read_add(VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z2n5;
wire VMR_L6D4_VMS_L6D4PHI3Z2n5_wr_en;
wire [5:0] VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2_number;
wire [10:0] VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2;
VMStubs #("Match") VMS_L6D4PHI3Z2n5(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z2n5),
.enable(VMR_L6D4_VMS_L6D4PHI3Z2n5_wr_en),
.number_out(VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2_number),
.read_add(VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2_read_add),
.data_out(VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z1;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1_read_add;
wire [12:0] VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1;
VMProjections  VMPROJ_L3L4_L6D4PHI4Z1(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z1),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z1_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1_number),
.read_add(VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI4Z1n3;
wire VMR_L6D4_VMS_L6D4PHI4Z1n3_wr_en;
wire [5:0] VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1_number;
wire [10:0] VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1_read_add;
wire [17:0] VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1;
VMStubs #("Match") VMS_L6D4PHI4Z1n3(
.data_in(VMR_L6D4_VMS_L6D4PHI4Z1n3),
.enable(VMR_L6D4_VMS_L6D4PHI4Z1n3_wr_en),
.number_out(VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1_number),
.read_add(VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1_read_add),
.data_out(VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z2;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2_read_add;
wire [12:0] VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2;
VMProjections  VMPROJ_L3L4_L6D4PHI4Z2(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z2),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z2_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2_number),
.read_add(VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI4Z2n3;
wire VMR_L6D4_VMS_L6D4PHI4Z2n3_wr_en;
wire [5:0] VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2_number;
wire [10:0] VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2_read_add;
wire [17:0] VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2;
VMStubs #("Match") VMS_L6D4PHI4Z2n3(
.data_in(VMR_L6D4_VMS_L6D4PHI4Z2n3),
.enable(VMR_L6D4_VMS_L6D4PHI4Z2n3_wr_en),
.number_out(VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2_number),
.read_add(VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2_read_add),
.data_out(VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z1;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1;
VMProjections  VMPROJ_L1L2_L3D3PHI1Z1(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z1),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z1_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1_number),
.read_add(VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z1n5;
wire VMR_L3D3_VMS_L3D3PHI1Z1n5_wr_en;
wire [5:0] VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1_number;
wire [10:0] VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1_read_add;
wire [17:0] VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1;
VMStubs #("Match") VMS_L3D3PHI1Z1n5(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z1n5),
.enable(VMR_L3D3_VMS_L3D3PHI1Z1n5_wr_en),
.number_out(VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1_number),
.read_add(VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1_read_add),
.data_out(VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z2;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2;
VMProjections  VMPROJ_L1L2_L3D3PHI1Z2(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z2),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z2_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2_number),
.read_add(VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z2n5;
wire VMR_L3D3_VMS_L3D3PHI1Z2n5_wr_en;
wire [5:0] VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2_number;
wire [10:0] VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2_read_add;
wire [17:0] VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2;
VMStubs #("Match") VMS_L3D3PHI1Z2n5(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z2n5),
.enable(VMR_L3D3_VMS_L3D3PHI1Z2n5_wr_en),
.number_out(VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2_number),
.read_add(VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2_read_add),
.data_out(VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z1;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1;
VMProjections  VMPROJ_L1L2_L3D3PHI2Z1(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z1),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z1_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1_number),
.read_add(VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z1n5;
wire VMR_L3D3_VMS_L3D3PHI2Z1n5_wr_en;
wire [5:0] VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1_number;
wire [10:0] VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1_read_add;
wire [17:0] VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1;
VMStubs #("Match") VMS_L3D3PHI2Z1n5(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z1n5),
.enable(VMR_L3D3_VMS_L3D3PHI2Z1n5_wr_en),
.number_out(VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1_number),
.read_add(VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1_read_add),
.data_out(VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z2;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2;
VMProjections  VMPROJ_L1L2_L3D3PHI2Z2(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z2),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z2_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2_number),
.read_add(VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z2n5;
wire VMR_L3D3_VMS_L3D3PHI2Z2n5_wr_en;
wire [5:0] VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2_number;
wire [10:0] VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2_read_add;
wire [17:0] VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2;
VMStubs #("Match") VMS_L3D3PHI2Z2n5(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z2n5),
.enable(VMR_L3D3_VMS_L3D3PHI2Z2n5_wr_en),
.number_out(VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2_number),
.read_add(VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2_read_add),
.data_out(VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z1;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1;
VMProjections  VMPROJ_L1L2_L3D3PHI3Z1(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z1),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z1_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1_number),
.read_add(VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z1n5;
wire VMR_L3D3_VMS_L3D3PHI3Z1n5_wr_en;
wire [5:0] VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1_number;
wire [10:0] VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1_read_add;
wire [17:0] VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1;
VMStubs #("Match") VMS_L3D3PHI3Z1n5(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z1n5),
.enable(VMR_L3D3_VMS_L3D3PHI3Z1n5_wr_en),
.number_out(VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1_number),
.read_add(VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1_read_add),
.data_out(VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z2;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2;
VMProjections  VMPROJ_L1L2_L3D3PHI3Z2(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z2),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z2_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2_number),
.read_add(VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z2n5;
wire VMR_L3D3_VMS_L3D3PHI3Z2n5_wr_en;
wire [5:0] VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2_number;
wire [10:0] VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2_read_add;
wire [17:0] VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2;
VMStubs #("Match") VMS_L3D3PHI3Z2n5(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z2n5),
.enable(VMR_L3D3_VMS_L3D3PHI3Z2n5_wr_en),
.number_out(VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2_number),
.read_add(VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2_read_add),
.data_out(VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z1;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1;
VMProjections  VMPROJ_L1L2_L3D4PHI1Z1(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z1),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z1_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1_number),
.read_add(VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z1n5;
wire VMR_L3D4_VMS_L3D4PHI1Z1n5_wr_en;
wire [5:0] VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1_number;
wire [10:0] VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1_read_add;
wire [17:0] VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1;
VMStubs #("Match") VMS_L3D4PHI1Z1n5(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z1n5),
.enable(VMR_L3D4_VMS_L3D4PHI1Z1n5_wr_en),
.number_out(VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1_number),
.read_add(VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1_read_add),
.data_out(VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z2;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2;
VMProjections  VMPROJ_L1L2_L3D4PHI1Z2(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z2),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z2_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2_number),
.read_add(VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z2n3;
wire VMR_L3D4_VMS_L3D4PHI1Z2n3_wr_en;
wire [5:0] VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2_number;
wire [10:0] VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2_read_add;
wire [17:0] VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2;
VMStubs #("Match") VMS_L3D4PHI1Z2n3(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z2n3),
.enable(VMR_L3D4_VMS_L3D4PHI1Z2n3_wr_en),
.number_out(VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2_number),
.read_add(VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2_read_add),
.data_out(VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z1;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1;
VMProjections  VMPROJ_L1L2_L3D4PHI2Z1(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z1),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z1_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1_number),
.read_add(VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z1n5;
wire VMR_L3D4_VMS_L3D4PHI2Z1n5_wr_en;
wire [5:0] VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1_number;
wire [10:0] VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1_read_add;
wire [17:0] VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1;
VMStubs #("Match") VMS_L3D4PHI2Z1n5(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z1n5),
.enable(VMR_L3D4_VMS_L3D4PHI2Z1n5_wr_en),
.number_out(VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1_number),
.read_add(VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1_read_add),
.data_out(VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z2;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2;
VMProjections  VMPROJ_L1L2_L3D4PHI2Z2(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z2),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z2_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2_number),
.read_add(VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z2n3;
wire VMR_L3D4_VMS_L3D4PHI2Z2n3_wr_en;
wire [5:0] VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2_number;
wire [10:0] VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2_read_add;
wire [17:0] VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2;
VMStubs #("Match") VMS_L3D4PHI2Z2n3(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z2n3),
.enable(VMR_L3D4_VMS_L3D4PHI2Z2n3_wr_en),
.number_out(VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2_number),
.read_add(VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2_read_add),
.data_out(VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z1;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1;
VMProjections  VMPROJ_L1L2_L3D4PHI3Z1(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z1),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z1_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1_number),
.read_add(VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z1n5;
wire VMR_L3D4_VMS_L3D4PHI3Z1n5_wr_en;
wire [5:0] VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1_number;
wire [10:0] VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1_read_add;
wire [17:0] VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1;
VMStubs #("Match") VMS_L3D4PHI3Z1n5(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z1n5),
.enable(VMR_L3D4_VMS_L3D4PHI3Z1n5_wr_en),
.number_out(VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1_number),
.read_add(VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1_read_add),
.data_out(VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z2;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2;
VMProjections  VMPROJ_L1L2_L3D4PHI3Z2(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z2),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z2_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2_number),
.read_add(VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z2n3;
wire VMR_L3D4_VMS_L3D4PHI3Z2n3_wr_en;
wire [5:0] VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2_number;
wire [10:0] VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2_read_add;
wire [17:0] VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2;
VMStubs #("Match") VMS_L3D4PHI3Z2n3(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z2n3),
.enable(VMR_L3D4_VMS_L3D4PHI3Z2n3_wr_en),
.number_out(VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2_number),
.read_add(VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2_read_add),
.data_out(VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z1;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1;
VMProjections  VMPROJ_L1L2_L4D3PHI1Z1(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z1),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z1_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1_number),
.read_add(VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI1Z1n2;
wire VMR_L4D3_VMS_L4D3PHI1Z1n2_wr_en;
wire [5:0] VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1_number;
wire [10:0] VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1_read_add;
wire [17:0] VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1;
VMStubs #("Match") VMS_L4D3PHI1Z1n2(
.data_in(VMR_L4D3_VMS_L4D3PHI1Z1n2),
.enable(VMR_L4D3_VMS_L4D3PHI1Z1n2_wr_en),
.number_out(VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1_number),
.read_add(VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1_read_add),
.data_out(VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z2;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2;
VMProjections  VMPROJ_L1L2_L4D3PHI1Z2(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z2),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z2_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2_number),
.read_add(VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI1Z2n3;
wire VMR_L4D3_VMS_L4D3PHI1Z2n3_wr_en;
wire [5:0] VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2_number;
wire [10:0] VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2_read_add;
wire [17:0] VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2;
VMStubs #("Match") VMS_L4D3PHI1Z2n3(
.data_in(VMR_L4D3_VMS_L4D3PHI1Z2n3),
.enable(VMR_L4D3_VMS_L4D3PHI1Z2n3_wr_en),
.number_out(VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2_number),
.read_add(VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2_read_add),
.data_out(VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z1;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1;
VMProjections  VMPROJ_L1L2_L4D3PHI2Z1(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z1),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z1_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1_number),
.read_add(VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z1n3;
wire VMR_L4D3_VMS_L4D3PHI2Z1n3_wr_en;
wire [5:0] VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1_number;
wire [10:0] VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1_read_add;
wire [17:0] VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1;
VMStubs #("Match") VMS_L4D3PHI2Z1n3(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z1n3),
.enable(VMR_L4D3_VMS_L4D3PHI2Z1n3_wr_en),
.number_out(VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1_number),
.read_add(VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1_read_add),
.data_out(VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z2;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2;
VMProjections  VMPROJ_L1L2_L4D3PHI2Z2(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z2),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z2_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2_number),
.read_add(VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z2n5;
wire VMR_L4D3_VMS_L4D3PHI2Z2n5_wr_en;
wire [5:0] VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2_number;
wire [10:0] VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2;
VMStubs #("Match") VMS_L4D3PHI2Z2n5(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z2n5),
.enable(VMR_L4D3_VMS_L4D3PHI2Z2n5_wr_en),
.number_out(VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2_number),
.read_add(VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2_read_add),
.data_out(VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z1;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1;
VMProjections  VMPROJ_L1L2_L4D3PHI3Z1(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z1),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z1_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1_number),
.read_add(VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z1n3;
wire VMR_L4D3_VMS_L4D3PHI3Z1n3_wr_en;
wire [5:0] VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1_number;
wire [10:0] VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1_read_add;
wire [17:0] VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1;
VMStubs #("Match") VMS_L4D3PHI3Z1n3(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z1n3),
.enable(VMR_L4D3_VMS_L4D3PHI3Z1n3_wr_en),
.number_out(VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1_number),
.read_add(VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1_read_add),
.data_out(VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z2;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2;
VMProjections  VMPROJ_L1L2_L4D3PHI3Z2(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z2),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z2_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2_number),
.read_add(VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z2n5;
wire VMR_L4D3_VMS_L4D3PHI3Z2n5_wr_en;
wire [5:0] VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2_number;
wire [10:0] VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2;
VMStubs #("Match") VMS_L4D3PHI3Z2n5(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z2n5),
.enable(VMR_L4D3_VMS_L4D3PHI3Z2n5_wr_en),
.number_out(VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2_number),
.read_add(VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2_read_add),
.data_out(VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z1;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1_read_add;
wire [12:0] VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1;
VMProjections  VMPROJ_L1L2_L4D3PHI4Z1(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z1),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z1_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1_number),
.read_add(VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI4Z1n2;
wire VMR_L4D3_VMS_L4D3PHI4Z1n2_wr_en;
wire [5:0] VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1_number;
wire [10:0] VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1_read_add;
wire [17:0] VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1;
VMStubs #("Match") VMS_L4D3PHI4Z1n2(
.data_in(VMR_L4D3_VMS_L4D3PHI4Z1n2),
.enable(VMR_L4D3_VMS_L4D3PHI4Z1n2_wr_en),
.number_out(VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1_number),
.read_add(VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1_read_add),
.data_out(VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z2;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2_read_add;
wire [12:0] VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2;
VMProjections  VMPROJ_L1L2_L4D3PHI4Z2(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z2),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z2_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2_number),
.read_add(VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI4Z2n3;
wire VMR_L4D3_VMS_L4D3PHI4Z2n3_wr_en;
wire [5:0] VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2_number;
wire [10:0] VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2_read_add;
wire [17:0] VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2;
VMStubs #("Match") VMS_L4D3PHI4Z2n3(
.data_in(VMR_L4D3_VMS_L4D3PHI4Z2n3),
.enable(VMR_L4D3_VMS_L4D3PHI4Z2n3_wr_en),
.number_out(VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2_number),
.read_add(VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2_read_add),
.data_out(VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z1;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1;
VMProjections  VMPROJ_L1L2_L4D4PHI1Z1(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z1),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z1_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1_number),
.read_add(VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI1Z1n3;
wire VMR_L4D4_VMS_L4D4PHI1Z1n3_wr_en;
wire [5:0] VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1_number;
wire [10:0] VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1_read_add;
wire [17:0] VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1;
VMStubs #("Match") VMS_L4D4PHI1Z1n3(
.data_in(VMR_L4D4_VMS_L4D4PHI1Z1n3),
.enable(VMR_L4D4_VMS_L4D4PHI1Z1n3_wr_en),
.number_out(VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1_number),
.read_add(VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1_read_add),
.data_out(VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z2;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2;
VMProjections  VMPROJ_L1L2_L4D4PHI1Z2(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z2),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z2_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2_number),
.read_add(VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI1Z2n3;
wire VMR_L4D4_VMS_L4D4PHI1Z2n3_wr_en;
wire [5:0] VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2_number;
wire [10:0] VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2_read_add;
wire [17:0] VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2;
VMStubs #("Match") VMS_L4D4PHI1Z2n3(
.data_in(VMR_L4D4_VMS_L4D4PHI1Z2n3),
.enable(VMR_L4D4_VMS_L4D4PHI1Z2n3_wr_en),
.number_out(VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2_number),
.read_add(VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2_read_add),
.data_out(VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z1;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1;
VMProjections  VMPROJ_L1L2_L4D4PHI2Z1(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z1),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z1_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1_number),
.read_add(VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z1n5;
wire VMR_L4D4_VMS_L4D4PHI2Z1n5_wr_en;
wire [5:0] VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1_number;
wire [10:0] VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1;
VMStubs #("Match") VMS_L4D4PHI2Z1n5(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z1n5),
.enable(VMR_L4D4_VMS_L4D4PHI2Z1n5_wr_en),
.number_out(VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1_number),
.read_add(VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1_read_add),
.data_out(VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z2;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2;
VMProjections  VMPROJ_L1L2_L4D4PHI2Z2(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z2),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z2_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2_number),
.read_add(VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z2n5;
wire VMR_L4D4_VMS_L4D4PHI2Z2n5_wr_en;
wire [5:0] VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2_number;
wire [10:0] VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2;
VMStubs #("Match") VMS_L4D4PHI2Z2n5(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z2n5),
.enable(VMR_L4D4_VMS_L4D4PHI2Z2n5_wr_en),
.number_out(VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2_number),
.read_add(VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2_read_add),
.data_out(VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z1;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1;
VMProjections  VMPROJ_L1L2_L4D4PHI3Z1(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z1),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z1_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1_number),
.read_add(VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z1n5;
wire VMR_L4D4_VMS_L4D4PHI3Z1n5_wr_en;
wire [5:0] VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1_number;
wire [10:0] VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1;
VMStubs #("Match") VMS_L4D4PHI3Z1n5(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z1n5),
.enable(VMR_L4D4_VMS_L4D4PHI3Z1n5_wr_en),
.number_out(VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1_number),
.read_add(VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1_read_add),
.data_out(VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z2;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2;
VMProjections  VMPROJ_L1L2_L4D4PHI3Z2(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z2),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z2_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2_number),
.read_add(VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z2n5;
wire VMR_L4D4_VMS_L4D4PHI3Z2n5_wr_en;
wire [5:0] VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2_number;
wire [10:0] VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2;
VMStubs #("Match") VMS_L4D4PHI3Z2n5(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z2n5),
.enable(VMR_L4D4_VMS_L4D4PHI3Z2n5_wr_en),
.number_out(VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2_number),
.read_add(VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2_read_add),
.data_out(VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z1;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1_read_add;
wire [12:0] VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1;
VMProjections  VMPROJ_L1L2_L4D4PHI4Z1(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z1),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z1_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1_number),
.read_add(VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI4Z1n3;
wire VMR_L4D4_VMS_L4D4PHI4Z1n3_wr_en;
wire [5:0] VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1_number;
wire [10:0] VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1_read_add;
wire [17:0] VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1;
VMStubs #("Match") VMS_L4D4PHI4Z1n3(
.data_in(VMR_L4D4_VMS_L4D4PHI4Z1n3),
.enable(VMR_L4D4_VMS_L4D4PHI4Z1n3_wr_en),
.number_out(VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1_number),
.read_add(VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1_read_add),
.data_out(VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z2;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2_read_add;
wire [12:0] VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2;
VMProjections  VMPROJ_L1L2_L4D4PHI4Z2(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z2),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z2_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2_number),
.read_add(VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI4Z2n3;
wire VMR_L4D4_VMS_L4D4PHI4Z2n3_wr_en;
wire [5:0] VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2_number;
wire [10:0] VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2_read_add;
wire [17:0] VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2;
VMStubs #("Match") VMS_L4D4PHI4Z2n3(
.data_in(VMR_L4D4_VMS_L4D4PHI4Z2n3),
.enable(VMR_L4D4_VMS_L4D4PHI4Z2n3_wr_en),
.number_out(VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2_number),
.read_add(VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2_read_add),
.data_out(VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z1;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1;
VMProjections  VMPROJ_L1L2_L5D3PHI1Z1(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z1),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z1_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1_number),
.read_add(VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z1n6;
wire VMR_L5D3_VMS_L5D3PHI1Z1n6_wr_en;
wire [5:0] VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1_number;
wire [10:0] VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1_read_add;
wire [17:0] VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1;
VMStubs #("Match") VMS_L5D3PHI1Z1n6(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z1n6),
.enable(VMR_L5D3_VMS_L5D3PHI1Z1n6_wr_en),
.number_out(VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1_number),
.read_add(VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1_read_add),
.data_out(VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z2;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2;
VMProjections  VMPROJ_L1L2_L5D3PHI1Z2(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z2),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z2_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2_number),
.read_add(VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI1Z2n6;
wire VMR_L5D3_VMS_L5D3PHI1Z2n6_wr_en;
wire [5:0] VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2_number;
wire [10:0] VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2_read_add;
wire [17:0] VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2;
VMStubs #("Match") VMS_L5D3PHI1Z2n6(
.data_in(VMR_L5D3_VMS_L5D3PHI1Z2n6),
.enable(VMR_L5D3_VMS_L5D3PHI1Z2n6_wr_en),
.number_out(VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2_number),
.read_add(VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2_read_add),
.data_out(VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z1;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1;
VMProjections  VMPROJ_L1L2_L5D3PHI2Z1(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z1),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z1_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1_number),
.read_add(VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z1n6;
wire VMR_L5D3_VMS_L5D3PHI2Z1n6_wr_en;
wire [5:0] VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1_number;
wire [10:0] VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1_read_add;
wire [17:0] VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1;
VMStubs #("Match") VMS_L5D3PHI2Z1n6(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z1n6),
.enable(VMR_L5D3_VMS_L5D3PHI2Z1n6_wr_en),
.number_out(VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1_number),
.read_add(VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1_read_add),
.data_out(VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z2;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2;
VMProjections  VMPROJ_L1L2_L5D3PHI2Z2(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z2),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z2_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2_number),
.read_add(VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI2Z2n6;
wire VMR_L5D3_VMS_L5D3PHI2Z2n6_wr_en;
wire [5:0] VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2_number;
wire [10:0] VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2_read_add;
wire [17:0] VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2;
VMStubs #("Match") VMS_L5D3PHI2Z2n6(
.data_in(VMR_L5D3_VMS_L5D3PHI2Z2n6),
.enable(VMR_L5D3_VMS_L5D3PHI2Z2n6_wr_en),
.number_out(VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2_number),
.read_add(VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2_read_add),
.data_out(VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z1;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1;
VMProjections  VMPROJ_L1L2_L5D3PHI3Z1(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z1),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z1_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1_number),
.read_add(VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z1n6;
wire VMR_L5D3_VMS_L5D3PHI3Z1n6_wr_en;
wire [5:0] VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1_number;
wire [10:0] VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1_read_add;
wire [17:0] VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1;
VMStubs #("Match") VMS_L5D3PHI3Z1n6(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z1n6),
.enable(VMR_L5D3_VMS_L5D3PHI3Z1n6_wr_en),
.number_out(VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1_number),
.read_add(VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1_read_add),
.data_out(VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z2;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2;
VMProjections  VMPROJ_L1L2_L5D3PHI3Z2(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z2),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z2_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2_number),
.read_add(VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D3_VMS_L5D3PHI3Z2n6;
wire VMR_L5D3_VMS_L5D3PHI3Z2n6_wr_en;
wire [5:0] VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2_number;
wire [10:0] VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2_read_add;
wire [17:0] VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2;
VMStubs #("Match") VMS_L5D3PHI3Z2n6(
.data_in(VMR_L5D3_VMS_L5D3PHI3Z2n6),
.enable(VMR_L5D3_VMS_L5D3PHI3Z2n6_wr_en),
.number_out(VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2_number),
.read_add(VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2_read_add),
.data_out(VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z1;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1;
VMProjections  VMPROJ_L1L2_L5D4PHI1Z1(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z1),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z1_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1_number),
.read_add(VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z1n6;
wire VMR_L5D4_VMS_L5D4PHI1Z1n6_wr_en;
wire [5:0] VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1_number;
wire [10:0] VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1_read_add;
wire [17:0] VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1;
VMStubs #("Match") VMS_L5D4PHI1Z1n6(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z1n6),
.enable(VMR_L5D4_VMS_L5D4PHI1Z1n6_wr_en),
.number_out(VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1_number),
.read_add(VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1_read_add),
.data_out(VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z2;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2;
VMProjections  VMPROJ_L1L2_L5D4PHI1Z2(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z2),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z2_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2_number),
.read_add(VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI1Z2n4;
wire VMR_L5D4_VMS_L5D4PHI1Z2n4_wr_en;
wire [5:0] VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2_number;
wire [10:0] VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2_read_add;
wire [17:0] VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2;
VMStubs #("Match") VMS_L5D4PHI1Z2n4(
.data_in(VMR_L5D4_VMS_L5D4PHI1Z2n4),
.enable(VMR_L5D4_VMS_L5D4PHI1Z2n4_wr_en),
.number_out(VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2_number),
.read_add(VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2_read_add),
.data_out(VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z1;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1;
VMProjections  VMPROJ_L1L2_L5D4PHI2Z1(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z1),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z1_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1_number),
.read_add(VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z1n6;
wire VMR_L5D4_VMS_L5D4PHI2Z1n6_wr_en;
wire [5:0] VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1_number;
wire [10:0] VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1_read_add;
wire [17:0] VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1;
VMStubs #("Match") VMS_L5D4PHI2Z1n6(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z1n6),
.enable(VMR_L5D4_VMS_L5D4PHI2Z1n6_wr_en),
.number_out(VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1_number),
.read_add(VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1_read_add),
.data_out(VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z2;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2;
VMProjections  VMPROJ_L1L2_L5D4PHI2Z2(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z2),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z2_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2_number),
.read_add(VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI2Z2n4;
wire VMR_L5D4_VMS_L5D4PHI2Z2n4_wr_en;
wire [5:0] VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2_number;
wire [10:0] VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2_read_add;
wire [17:0] VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2;
VMStubs #("Match") VMS_L5D4PHI2Z2n4(
.data_in(VMR_L5D4_VMS_L5D4PHI2Z2n4),
.enable(VMR_L5D4_VMS_L5D4PHI2Z2n4_wr_en),
.number_out(VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2_number),
.read_add(VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2_read_add),
.data_out(VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z1;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1;
VMProjections  VMPROJ_L1L2_L5D4PHI3Z1(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z1),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z1_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1_number),
.read_add(VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z1n6;
wire VMR_L5D4_VMS_L5D4PHI3Z1n6_wr_en;
wire [5:0] VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1_number;
wire [10:0] VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1_read_add;
wire [17:0] VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1;
VMStubs #("Match") VMS_L5D4PHI3Z1n6(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z1n6),
.enable(VMR_L5D4_VMS_L5D4PHI3Z1n6_wr_en),
.number_out(VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1_number),
.read_add(VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1_read_add),
.data_out(VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z2;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2;
VMProjections  VMPROJ_L1L2_L5D4PHI3Z2(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z2),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z2_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2_number),
.read_add(VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L5D4_VMS_L5D4PHI3Z2n4;
wire VMR_L5D4_VMS_L5D4PHI3Z2n4_wr_en;
wire [5:0] VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2_number;
wire [10:0] VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2_read_add;
wire [17:0] VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2;
VMStubs #("Match") VMS_L5D4PHI3Z2n4(
.data_in(VMR_L5D4_VMS_L5D4PHI3Z2n4),
.enable(VMR_L5D4_VMS_L5D4PHI3Z2n4_wr_en),
.number_out(VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2_number),
.read_add(VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2_read_add),
.data_out(VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z1;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1;
VMProjections  VMPROJ_L1L2_L6D3PHI1Z1(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z1),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z1_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1_number),
.read_add(VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI1Z1n3;
wire VMR_L6D3_VMS_L6D3PHI1Z1n3_wr_en;
wire [5:0] VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1_number;
wire [10:0] VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1_read_add;
wire [17:0] VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1;
VMStubs #("Match") VMS_L6D3PHI1Z1n3(
.data_in(VMR_L6D3_VMS_L6D3PHI1Z1n3),
.enable(VMR_L6D3_VMS_L6D3PHI1Z1n3_wr_en),
.number_out(VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1_number),
.read_add(VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1_read_add),
.data_out(VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z2;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2;
VMProjections  VMPROJ_L1L2_L6D3PHI1Z2(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z2),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z2_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2_number),
.read_add(VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI1Z2n4;
wire VMR_L6D3_VMS_L6D3PHI1Z2n4_wr_en;
wire [5:0] VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2_number;
wire [10:0] VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2_read_add;
wire [17:0] VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2;
VMStubs #("Match") VMS_L6D3PHI1Z2n4(
.data_in(VMR_L6D3_VMS_L6D3PHI1Z2n4),
.enable(VMR_L6D3_VMS_L6D3PHI1Z2n4_wr_en),
.number_out(VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2_number),
.read_add(VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2_read_add),
.data_out(VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z1;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1;
VMProjections  VMPROJ_L1L2_L6D3PHI2Z1(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z1),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z1_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1_number),
.read_add(VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z1n4;
wire VMR_L6D3_VMS_L6D3PHI2Z1n4_wr_en;
wire [5:0] VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1_number;
wire [10:0] VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1_read_add;
wire [17:0] VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1;
VMStubs #("Match") VMS_L6D3PHI2Z1n4(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z1n4),
.enable(VMR_L6D3_VMS_L6D3PHI2Z1n4_wr_en),
.number_out(VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1_number),
.read_add(VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1_read_add),
.data_out(VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z2;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2;
VMProjections  VMPROJ_L1L2_L6D3PHI2Z2(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z2),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z2_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2_number),
.read_add(VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI2Z2n6;
wire VMR_L6D3_VMS_L6D3PHI2Z2n6_wr_en;
wire [5:0] VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2_number;
wire [10:0] VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2_read_add;
wire [17:0] VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2;
VMStubs #("Match") VMS_L6D3PHI2Z2n6(
.data_in(VMR_L6D3_VMS_L6D3PHI2Z2n6),
.enable(VMR_L6D3_VMS_L6D3PHI2Z2n6_wr_en),
.number_out(VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2_number),
.read_add(VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2_read_add),
.data_out(VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z1;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1;
VMProjections  VMPROJ_L1L2_L6D3PHI3Z1(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z1),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z1_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1_number),
.read_add(VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z1n4;
wire VMR_L6D3_VMS_L6D3PHI3Z1n4_wr_en;
wire [5:0] VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1_number;
wire [10:0] VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1_read_add;
wire [17:0] VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1;
VMStubs #("Match") VMS_L6D3PHI3Z1n4(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z1n4),
.enable(VMR_L6D3_VMS_L6D3PHI3Z1n4_wr_en),
.number_out(VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1_number),
.read_add(VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1_read_add),
.data_out(VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z2;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2;
VMProjections  VMPROJ_L1L2_L6D3PHI3Z2(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z2),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z2_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2_number),
.read_add(VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI3Z2n6;
wire VMR_L6D3_VMS_L6D3PHI3Z2n6_wr_en;
wire [5:0] VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2_number;
wire [10:0] VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2_read_add;
wire [17:0] VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2;
VMStubs #("Match") VMS_L6D3PHI3Z2n6(
.data_in(VMR_L6D3_VMS_L6D3PHI3Z2n6),
.enable(VMR_L6D3_VMS_L6D3PHI3Z2n6_wr_en),
.number_out(VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2_number),
.read_add(VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2_read_add),
.data_out(VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z1;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1_read_add;
wire [12:0] VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1;
VMProjections  VMPROJ_L1L2_L6D3PHI4Z1(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z1),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z1_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1_number),
.read_add(VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI4Z1n3;
wire VMR_L6D3_VMS_L6D3PHI4Z1n3_wr_en;
wire [5:0] VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1_number;
wire [10:0] VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1_read_add;
wire [17:0] VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1;
VMStubs #("Match") VMS_L6D3PHI4Z1n3(
.data_in(VMR_L6D3_VMS_L6D3PHI4Z1n3),
.enable(VMR_L6D3_VMS_L6D3PHI4Z1n3_wr_en),
.number_out(VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1_number),
.read_add(VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1_read_add),
.data_out(VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z2;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2_read_add;
wire [12:0] VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2;
VMProjections  VMPROJ_L1L2_L6D3PHI4Z2(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z2),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z2_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2_number),
.read_add(VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D3_VMS_L6D3PHI4Z2n4;
wire VMR_L6D3_VMS_L6D3PHI4Z2n4_wr_en;
wire [5:0] VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2_number;
wire [10:0] VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2_read_add;
wire [17:0] VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2;
VMStubs #("Match") VMS_L6D3PHI4Z2n4(
.data_in(VMR_L6D3_VMS_L6D3PHI4Z2n4),
.enable(VMR_L6D3_VMS_L6D3PHI4Z2n4_wr_en),
.number_out(VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2_number),
.read_add(VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2_read_add),
.data_out(VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z1;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1;
VMProjections  VMPROJ_L1L2_L6D4PHI1Z1(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z1),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z1_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1_number),
.read_add(VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI1Z1n4;
wire VMR_L6D4_VMS_L6D4PHI1Z1n4_wr_en;
wire [5:0] VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1_number;
wire [10:0] VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1_read_add;
wire [17:0] VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1;
VMStubs #("Match") VMS_L6D4PHI1Z1n4(
.data_in(VMR_L6D4_VMS_L6D4PHI1Z1n4),
.enable(VMR_L6D4_VMS_L6D4PHI1Z1n4_wr_en),
.number_out(VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1_number),
.read_add(VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1_read_add),
.data_out(VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z2;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2;
VMProjections  VMPROJ_L1L2_L6D4PHI1Z2(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z2),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z2_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2_number),
.read_add(VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI1Z2n4;
wire VMR_L6D4_VMS_L6D4PHI1Z2n4_wr_en;
wire [5:0] VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2_number;
wire [10:0] VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2_read_add;
wire [17:0] VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2;
VMStubs #("Match") VMS_L6D4PHI1Z2n4(
.data_in(VMR_L6D4_VMS_L6D4PHI1Z2n4),
.enable(VMR_L6D4_VMS_L6D4PHI1Z2n4_wr_en),
.number_out(VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2_number),
.read_add(VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2_read_add),
.data_out(VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z1;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1;
VMProjections  VMPROJ_L1L2_L6D4PHI2Z1(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z1),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z1_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1_number),
.read_add(VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z1n6;
wire VMR_L6D4_VMS_L6D4PHI2Z1n6_wr_en;
wire [5:0] VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1_number;
wire [10:0] VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1_read_add;
wire [17:0] VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1;
VMStubs #("Match") VMS_L6D4PHI2Z1n6(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z1n6),
.enable(VMR_L6D4_VMS_L6D4PHI2Z1n6_wr_en),
.number_out(VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1_number),
.read_add(VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1_read_add),
.data_out(VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z2;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2;
VMProjections  VMPROJ_L1L2_L6D4PHI2Z2(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z2),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z2_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2_number),
.read_add(VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI2Z2n6;
wire VMR_L6D4_VMS_L6D4PHI2Z2n6_wr_en;
wire [5:0] VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2_number;
wire [10:0] VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2_read_add;
wire [17:0] VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2;
VMStubs #("Match") VMS_L6D4PHI2Z2n6(
.data_in(VMR_L6D4_VMS_L6D4PHI2Z2n6),
.enable(VMR_L6D4_VMS_L6D4PHI2Z2n6_wr_en),
.number_out(VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2_number),
.read_add(VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2_read_add),
.data_out(VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z1;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1;
VMProjections  VMPROJ_L1L2_L6D4PHI3Z1(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z1),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z1_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1_number),
.read_add(VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z1n6;
wire VMR_L6D4_VMS_L6D4PHI3Z1n6_wr_en;
wire [5:0] VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1_number;
wire [10:0] VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1_read_add;
wire [17:0] VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1;
VMStubs #("Match") VMS_L6D4PHI3Z1n6(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z1n6),
.enable(VMR_L6D4_VMS_L6D4PHI3Z1n6_wr_en),
.number_out(VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1_number),
.read_add(VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1_read_add),
.data_out(VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z2;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2;
VMProjections  VMPROJ_L1L2_L6D4PHI3Z2(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z2),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z2_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2_number),
.read_add(VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI3Z2n6;
wire VMR_L6D4_VMS_L6D4PHI3Z2n6_wr_en;
wire [5:0] VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2_number;
wire [10:0] VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2_read_add;
wire [17:0] VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2;
VMStubs #("Match") VMS_L6D4PHI3Z2n6(
.data_in(VMR_L6D4_VMS_L6D4PHI3Z2n6),
.enable(VMR_L6D4_VMS_L6D4PHI3Z2n6_wr_en),
.number_out(VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2_number),
.read_add(VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2_read_add),
.data_out(VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z1;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1_read_add;
wire [12:0] VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1;
VMProjections  VMPROJ_L1L2_L6D4PHI4Z1(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z1),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z1_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1_number),
.read_add(VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI4Z1n4;
wire VMR_L6D4_VMS_L6D4PHI4Z1n4_wr_en;
wire [5:0] VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1_number;
wire [10:0] VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1_read_add;
wire [17:0] VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1;
VMStubs #("Match") VMS_L6D4PHI4Z1n4(
.data_in(VMR_L6D4_VMS_L6D4PHI4Z1n4),
.enable(VMR_L6D4_VMS_L6D4PHI4Z1n4_wr_en),
.number_out(VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1_number),
.read_add(VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1_read_add),
.data_out(VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z2;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2_read_add;
wire [12:0] VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2;
VMProjections  VMPROJ_L1L2_L6D4PHI4Z2(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z2),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z2_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2_number),
.read_add(VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L6D4_VMS_L6D4PHI4Z2n4;
wire VMR_L6D4_VMS_L6D4PHI4Z2n4_wr_en;
wire [5:0] VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2_number;
wire [10:0] VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2_read_add;
wire [17:0] VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2;
VMStubs #("Match") VMS_L6D4PHI4Z2n4(
.data_in(VMR_L6D4_VMS_L6D4PHI4Z2n4),
.enable(VMR_L6D4_VMS_L6D4PHI4Z2n4_wr_en),
.number_out(VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2_number),
.read_add(VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2_read_add),
.data_out(VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z1;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1;
VMProjections  VMPROJ_L5L6_L1D3PHI1Z1(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z1),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z1_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1_number),
.read_add(VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z1n8;
wire VMR_L1D3_VMS_L1D3PHI1Z1n8_wr_en;
wire [5:0] VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1_number;
wire [10:0] VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1_read_add;
wire [17:0] VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1;
VMStubs #("Match") VMS_L1D3PHI1Z1n8(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z1n8),
.enable(VMR_L1D3_VMS_L1D3PHI1Z1n8_wr_en),
.number_out(VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1_number),
.read_add(VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1_read_add),
.data_out(VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z2;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2;
VMProjections  VMPROJ_L5L6_L1D3PHI1Z2(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z2),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z2_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2_number),
.read_add(VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI1Z2n8;
wire VMR_L1D3_VMS_L1D3PHI1Z2n8_wr_en;
wire [5:0] VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2_number;
wire [10:0] VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2_read_add;
wire [17:0] VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2;
VMStubs #("Match") VMS_L1D3PHI1Z2n8(
.data_in(VMR_L1D3_VMS_L1D3PHI1Z2n8),
.enable(VMR_L1D3_VMS_L1D3PHI1Z2n8_wr_en),
.number_out(VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2_number),
.read_add(VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2_read_add),
.data_out(VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z1;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1;
VMProjections  VMPROJ_L5L6_L1D3PHI2Z1(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z1),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z1_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1_number),
.read_add(VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z1n8;
wire VMR_L1D3_VMS_L1D3PHI2Z1n8_wr_en;
wire [5:0] VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1_number;
wire [10:0] VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1_read_add;
wire [17:0] VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1;
VMStubs #("Match") VMS_L1D3PHI2Z1n8(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z1n8),
.enable(VMR_L1D3_VMS_L1D3PHI2Z1n8_wr_en),
.number_out(VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1_number),
.read_add(VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1_read_add),
.data_out(VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z2;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2;
VMProjections  VMPROJ_L5L6_L1D3PHI2Z2(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z2),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z2_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2_number),
.read_add(VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI2Z2n8;
wire VMR_L1D3_VMS_L1D3PHI2Z2n8_wr_en;
wire [5:0] VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2_number;
wire [10:0] VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2_read_add;
wire [17:0] VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2;
VMStubs #("Match") VMS_L1D3PHI2Z2n8(
.data_in(VMR_L1D3_VMS_L1D3PHI2Z2n8),
.enable(VMR_L1D3_VMS_L1D3PHI2Z2n8_wr_en),
.number_out(VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2_number),
.read_add(VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2_read_add),
.data_out(VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z1;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1;
VMProjections  VMPROJ_L5L6_L1D3PHI3Z1(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z1),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z1_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1_number),
.read_add(VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z1n8;
wire VMR_L1D3_VMS_L1D3PHI3Z1n8_wr_en;
wire [5:0] VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1_number;
wire [10:0] VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1_read_add;
wire [17:0] VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1;
VMStubs #("Match") VMS_L1D3PHI3Z1n8(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z1n8),
.enable(VMR_L1D3_VMS_L1D3PHI3Z1n8_wr_en),
.number_out(VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1_number),
.read_add(VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1_read_add),
.data_out(VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z2;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2;
VMProjections  VMPROJ_L5L6_L1D3PHI3Z2(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z2),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z2_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2_number),
.read_add(VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D3_VMS_L1D3PHI3Z2n8;
wire VMR_L1D3_VMS_L1D3PHI3Z2n8_wr_en;
wire [5:0] VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2_number;
wire [10:0] VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2_read_add;
wire [17:0] VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2;
VMStubs #("Match") VMS_L1D3PHI3Z2n8(
.data_in(VMR_L1D3_VMS_L1D3PHI3Z2n8),
.enable(VMR_L1D3_VMS_L1D3PHI3Z2n8_wr_en),
.number_out(VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2_number),
.read_add(VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2_read_add),
.data_out(VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z1;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1;
VMProjections  VMPROJ_L5L6_L1D4PHI1Z1(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z1),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z1_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1_number),
.read_add(VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI1Z1n4;
wire VMR_L1D4_VMS_L1D4PHI1Z1n4_wr_en;
wire [5:0] VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1_number;
wire [10:0] VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1_read_add;
wire [17:0] VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1;
VMStubs #("Match") VMS_L1D4PHI1Z1n4(
.data_in(VMR_L1D4_VMS_L1D4PHI1Z1n4),
.enable(VMR_L1D4_VMS_L1D4PHI1Z1n4_wr_en),
.number_out(VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1_number),
.read_add(VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1_read_add),
.data_out(VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z2;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2;
VMProjections  VMPROJ_L5L6_L1D4PHI1Z2(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z2),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z2_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2_number),
.read_add(VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI1Z2n2;
wire VMR_L1D4_VMS_L1D4PHI1Z2n2_wr_en;
wire [5:0] VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2_number;
wire [10:0] VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2_read_add;
wire [17:0] VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2;
VMStubs #("Match") VMS_L1D4PHI1Z2n2(
.data_in(VMR_L1D4_VMS_L1D4PHI1Z2n2),
.enable(VMR_L1D4_VMS_L1D4PHI1Z2n2_wr_en),
.number_out(VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2_number),
.read_add(VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2_read_add),
.data_out(VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z1;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1;
VMProjections  VMPROJ_L5L6_L1D4PHI2Z1(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z1),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z1_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1_number),
.read_add(VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI2Z1n4;
wire VMR_L1D4_VMS_L1D4PHI2Z1n4_wr_en;
wire [5:0] VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1_number;
wire [10:0] VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1_read_add;
wire [17:0] VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1;
VMStubs #("Match") VMS_L1D4PHI2Z1n4(
.data_in(VMR_L1D4_VMS_L1D4PHI2Z1n4),
.enable(VMR_L1D4_VMS_L1D4PHI2Z1n4_wr_en),
.number_out(VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1_number),
.read_add(VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1_read_add),
.data_out(VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z2;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2;
VMProjections  VMPROJ_L5L6_L1D4PHI2Z2(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z2),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z2_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2_number),
.read_add(VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI2Z2n2;
wire VMR_L1D4_VMS_L1D4PHI2Z2n2_wr_en;
wire [5:0] VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2_number;
wire [10:0] VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2_read_add;
wire [17:0] VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2;
VMStubs #("Match") VMS_L1D4PHI2Z2n2(
.data_in(VMR_L1D4_VMS_L1D4PHI2Z2n2),
.enable(VMR_L1D4_VMS_L1D4PHI2Z2n2_wr_en),
.number_out(VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2_number),
.read_add(VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2_read_add),
.data_out(VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z1;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1;
VMProjections  VMPROJ_L5L6_L1D4PHI3Z1(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z1),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z1_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1_number),
.read_add(VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI3Z1n4;
wire VMR_L1D4_VMS_L1D4PHI3Z1n4_wr_en;
wire [5:0] VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1_number;
wire [10:0] VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1_read_add;
wire [17:0] VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1;
VMStubs #("Match") VMS_L1D4PHI3Z1n4(
.data_in(VMR_L1D4_VMS_L1D4PHI3Z1n4),
.enable(VMR_L1D4_VMS_L1D4PHI3Z1n4_wr_en),
.number_out(VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1_number),
.read_add(VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1_read_add),
.data_out(VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z2;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2;
VMProjections  VMPROJ_L5L6_L1D4PHI3Z2(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z2),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z2_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2_number),
.read_add(VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L1D4_VMS_L1D4PHI3Z2n2;
wire VMR_L1D4_VMS_L1D4PHI3Z2n2_wr_en;
wire [5:0] VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2_number;
wire [10:0] VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2_read_add;
wire [17:0] VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2;
VMStubs #("Match") VMS_L1D4PHI3Z2n2(
.data_in(VMR_L1D4_VMS_L1D4PHI3Z2n2),
.enable(VMR_L1D4_VMS_L1D4PHI3Z2n2_wr_en),
.number_out(VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2_number),
.read_add(VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2_read_add),
.data_out(VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z1;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1;
VMProjections  VMPROJ_L5L6_L2D3PHI1Z1(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z1),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z1_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1_number),
.read_add(VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI1Z1n3;
wire VMR_L2D3_VMS_L2D3PHI1Z1n3_wr_en;
wire [5:0] VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1_number;
wire [10:0] VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1_read_add;
wire [17:0] VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1;
VMStubs #("Match") VMS_L2D3PHI1Z1n3(
.data_in(VMR_L2D3_VMS_L2D3PHI1Z1n3),
.enable(VMR_L2D3_VMS_L2D3PHI1Z1n3_wr_en),
.number_out(VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1_number),
.read_add(VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1_read_add),
.data_out(VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z2;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2;
VMProjections  VMPROJ_L5L6_L2D3PHI1Z2(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z2),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z2_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2_number),
.read_add(VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI1Z2n4;
wire VMR_L2D3_VMS_L2D3PHI1Z2n4_wr_en;
wire [5:0] VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2_number;
wire [10:0] VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2_read_add;
wire [17:0] VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2;
VMStubs #("Match") VMS_L2D3PHI1Z2n4(
.data_in(VMR_L2D3_VMS_L2D3PHI1Z2n4),
.enable(VMR_L2D3_VMS_L2D3PHI1Z2n4_wr_en),
.number_out(VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2_number),
.read_add(VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2_read_add),
.data_out(VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z1;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1;
VMProjections  VMPROJ_L5L6_L2D3PHI2Z1(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z1),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z1_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1_number),
.read_add(VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z1n4;
wire VMR_L2D3_VMS_L2D3PHI2Z1n4_wr_en;
wire [5:0] VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1_number;
wire [10:0] VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1_read_add;
wire [17:0] VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1;
VMStubs #("Match") VMS_L2D3PHI2Z1n4(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z1n4),
.enable(VMR_L2D3_VMS_L2D3PHI2Z1n4_wr_en),
.number_out(VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1_number),
.read_add(VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1_read_add),
.data_out(VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z2;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2;
VMProjections  VMPROJ_L5L6_L2D3PHI2Z2(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z2),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z2_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2_number),
.read_add(VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI2Z2n6;
wire VMR_L2D3_VMS_L2D3PHI2Z2n6_wr_en;
wire [5:0] VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2_number;
wire [10:0] VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2_read_add;
wire [17:0] VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2;
VMStubs #("Match") VMS_L2D3PHI2Z2n6(
.data_in(VMR_L2D3_VMS_L2D3PHI2Z2n6),
.enable(VMR_L2D3_VMS_L2D3PHI2Z2n6_wr_en),
.number_out(VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2_number),
.read_add(VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2_read_add),
.data_out(VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z1;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1;
VMProjections  VMPROJ_L5L6_L2D3PHI3Z1(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z1),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z1_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1_number),
.read_add(VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z1n4;
wire VMR_L2D3_VMS_L2D3PHI3Z1n4_wr_en;
wire [5:0] VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1_number;
wire [10:0] VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1_read_add;
wire [17:0] VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1;
VMStubs #("Match") VMS_L2D3PHI3Z1n4(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z1n4),
.enable(VMR_L2D3_VMS_L2D3PHI3Z1n4_wr_en),
.number_out(VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1_number),
.read_add(VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1_read_add),
.data_out(VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z2;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2;
VMProjections  VMPROJ_L5L6_L2D3PHI3Z2(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z2),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z2_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2_number),
.read_add(VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI3Z2n6;
wire VMR_L2D3_VMS_L2D3PHI3Z2n6_wr_en;
wire [5:0] VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2_number;
wire [10:0] VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2_read_add;
wire [17:0] VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2;
VMStubs #("Match") VMS_L2D3PHI3Z2n6(
.data_in(VMR_L2D3_VMS_L2D3PHI3Z2n6),
.enable(VMR_L2D3_VMS_L2D3PHI3Z2n6_wr_en),
.number_out(VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2_number),
.read_add(VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2_read_add),
.data_out(VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z1;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1_read_add;
wire [12:0] VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1;
VMProjections  VMPROJ_L5L6_L2D3PHI4Z1(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z1),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z1_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1_number),
.read_add(VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI4Z1n3;
wire VMR_L2D3_VMS_L2D3PHI4Z1n3_wr_en;
wire [5:0] VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1_number;
wire [10:0] VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1_read_add;
wire [17:0] VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1;
VMStubs #("Match") VMS_L2D3PHI4Z1n3(
.data_in(VMR_L2D3_VMS_L2D3PHI4Z1n3),
.enable(VMR_L2D3_VMS_L2D3PHI4Z1n3_wr_en),
.number_out(VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1_number),
.read_add(VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1_read_add),
.data_out(VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z2;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2_read_add;
wire [12:0] VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2;
VMProjections  VMPROJ_L5L6_L2D3PHI4Z2(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z2),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z2_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2_number),
.read_add(VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D3_VMS_L2D3PHI4Z2n4;
wire VMR_L2D3_VMS_L2D3PHI4Z2n4_wr_en;
wire [5:0] VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2_number;
wire [10:0] VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2_read_add;
wire [17:0] VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2;
VMStubs #("Match") VMS_L2D3PHI4Z2n4(
.data_in(VMR_L2D3_VMS_L2D3PHI4Z2n4),
.enable(VMR_L2D3_VMS_L2D3PHI4Z2n4_wr_en),
.number_out(VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2_number),
.read_add(VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2_read_add),
.data_out(VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z1;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1;
VMProjections  VMPROJ_L5L6_L2D4PHI1Z1(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z1),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z1_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1_number),
.read_add(VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI1Z1n4;
wire VMR_L2D4_VMS_L2D4PHI1Z1n4_wr_en;
wire [5:0] VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1_number;
wire [10:0] VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1_read_add;
wire [17:0] VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1;
VMStubs #("Match") VMS_L2D4PHI1Z1n4(
.data_in(VMR_L2D4_VMS_L2D4PHI1Z1n4),
.enable(VMR_L2D4_VMS_L2D4PHI1Z1n4_wr_en),
.number_out(VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1_number),
.read_add(VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1_read_add),
.data_out(VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z2;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2;
VMProjections  VMPROJ_L5L6_L2D4PHI1Z2(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z2),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z2_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2_number),
.read_add(VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI1Z2n4;
wire VMR_L2D4_VMS_L2D4PHI1Z2n4_wr_en;
wire [5:0] VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2_number;
wire [10:0] VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2_read_add;
wire [17:0] VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2;
VMStubs #("Match") VMS_L2D4PHI1Z2n4(
.data_in(VMR_L2D4_VMS_L2D4PHI1Z2n4),
.enable(VMR_L2D4_VMS_L2D4PHI1Z2n4_wr_en),
.number_out(VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2_number),
.read_add(VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2_read_add),
.data_out(VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z1;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1;
VMProjections  VMPROJ_L5L6_L2D4PHI2Z1(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z1),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z1_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1_number),
.read_add(VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z1n6;
wire VMR_L2D4_VMS_L2D4PHI2Z1n6_wr_en;
wire [5:0] VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1_number;
wire [10:0] VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1_read_add;
wire [17:0] VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1;
VMStubs #("Match") VMS_L2D4PHI2Z1n6(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z1n6),
.enable(VMR_L2D4_VMS_L2D4PHI2Z1n6_wr_en),
.number_out(VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1_number),
.read_add(VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1_read_add),
.data_out(VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z2;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2;
VMProjections  VMPROJ_L5L6_L2D4PHI2Z2(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z2),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z2_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2_number),
.read_add(VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI2Z2n6;
wire VMR_L2D4_VMS_L2D4PHI2Z2n6_wr_en;
wire [5:0] VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2_number;
wire [10:0] VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2_read_add;
wire [17:0] VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2;
VMStubs #("Match") VMS_L2D4PHI2Z2n6(
.data_in(VMR_L2D4_VMS_L2D4PHI2Z2n6),
.enable(VMR_L2D4_VMS_L2D4PHI2Z2n6_wr_en),
.number_out(VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2_number),
.read_add(VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2_read_add),
.data_out(VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z1;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1;
VMProjections  VMPROJ_L5L6_L2D4PHI3Z1(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z1),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z1_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1_number),
.read_add(VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z1n6;
wire VMR_L2D4_VMS_L2D4PHI3Z1n6_wr_en;
wire [5:0] VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1_number;
wire [10:0] VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1_read_add;
wire [17:0] VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1;
VMStubs #("Match") VMS_L2D4PHI3Z1n6(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z1n6),
.enable(VMR_L2D4_VMS_L2D4PHI3Z1n6_wr_en),
.number_out(VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1_number),
.read_add(VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1_read_add),
.data_out(VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z2;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2;
VMProjections  VMPROJ_L5L6_L2D4PHI3Z2(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z2),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z2_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2_number),
.read_add(VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI3Z2n6;
wire VMR_L2D4_VMS_L2D4PHI3Z2n6_wr_en;
wire [5:0] VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2_number;
wire [10:0] VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2_read_add;
wire [17:0] VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2;
VMStubs #("Match") VMS_L2D4PHI3Z2n6(
.data_in(VMR_L2D4_VMS_L2D4PHI3Z2n6),
.enable(VMR_L2D4_VMS_L2D4PHI3Z2n6_wr_en),
.number_out(VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2_number),
.read_add(VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2_read_add),
.data_out(VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z1;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1_read_add;
wire [12:0] VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1;
VMProjections  VMPROJ_L5L6_L2D4PHI4Z1(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z1),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z1_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1_number),
.read_add(VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI4Z1n4;
wire VMR_L2D4_VMS_L2D4PHI4Z1n4_wr_en;
wire [5:0] VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1_number;
wire [10:0] VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1_read_add;
wire [17:0] VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1;
VMStubs #("Match") VMS_L2D4PHI4Z1n4(
.data_in(VMR_L2D4_VMS_L2D4PHI4Z1n4),
.enable(VMR_L2D4_VMS_L2D4PHI4Z1n4_wr_en),
.number_out(VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1_number),
.read_add(VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1_read_add),
.data_out(VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z2;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2_read_add;
wire [12:0] VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2;
VMProjections  VMPROJ_L5L6_L2D4PHI4Z2(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z2),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z2_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2_number),
.read_add(VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L2D4_VMS_L2D4PHI4Z2n4;
wire VMR_L2D4_VMS_L2D4PHI4Z2n4_wr_en;
wire [5:0] VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2_number;
wire [10:0] VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2_read_add;
wire [17:0] VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2;
VMStubs #("Match") VMS_L2D4PHI4Z2n4(
.data_in(VMR_L2D4_VMS_L2D4PHI4Z2n4),
.enable(VMR_L2D4_VMS_L2D4PHI4Z2n4_wr_en),
.number_out(VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2_number),
.read_add(VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2_read_add),
.data_out(VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z1;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1;
VMProjections  VMPROJ_L5L6_L3D3PHI1Z1(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z1),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z1_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1_number),
.read_add(VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z1n6;
wire VMR_L3D3_VMS_L3D3PHI1Z1n6_wr_en;
wire [5:0] VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1_number;
wire [10:0] VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1_read_add;
wire [17:0] VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1;
VMStubs #("Match") VMS_L3D3PHI1Z1n6(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z1n6),
.enable(VMR_L3D3_VMS_L3D3PHI1Z1n6_wr_en),
.number_out(VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1_number),
.read_add(VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1_read_add),
.data_out(VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z2;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2;
VMProjections  VMPROJ_L5L6_L3D3PHI1Z2(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z2),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z2_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2_number),
.read_add(VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI1Z2n6;
wire VMR_L3D3_VMS_L3D3PHI1Z2n6_wr_en;
wire [5:0] VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2_number;
wire [10:0] VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2_read_add;
wire [17:0] VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2;
VMStubs #("Match") VMS_L3D3PHI1Z2n6(
.data_in(VMR_L3D3_VMS_L3D3PHI1Z2n6),
.enable(VMR_L3D3_VMS_L3D3PHI1Z2n6_wr_en),
.number_out(VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2_number),
.read_add(VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2_read_add),
.data_out(VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z1;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1;
VMProjections  VMPROJ_L5L6_L3D3PHI2Z1(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z1),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z1_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1_number),
.read_add(VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z1n6;
wire VMR_L3D3_VMS_L3D3PHI2Z1n6_wr_en;
wire [5:0] VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1_number;
wire [10:0] VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1_read_add;
wire [17:0] VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1;
VMStubs #("Match") VMS_L3D3PHI2Z1n6(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z1n6),
.enable(VMR_L3D3_VMS_L3D3PHI2Z1n6_wr_en),
.number_out(VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1_number),
.read_add(VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1_read_add),
.data_out(VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z2;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2;
VMProjections  VMPROJ_L5L6_L3D3PHI2Z2(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z2),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z2_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2_number),
.read_add(VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI2Z2n6;
wire VMR_L3D3_VMS_L3D3PHI2Z2n6_wr_en;
wire [5:0] VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2_number;
wire [10:0] VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2_read_add;
wire [17:0] VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2;
VMStubs #("Match") VMS_L3D3PHI2Z2n6(
.data_in(VMR_L3D3_VMS_L3D3PHI2Z2n6),
.enable(VMR_L3D3_VMS_L3D3PHI2Z2n6_wr_en),
.number_out(VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2_number),
.read_add(VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2_read_add),
.data_out(VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z1;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1;
VMProjections  VMPROJ_L5L6_L3D3PHI3Z1(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z1),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z1_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1_number),
.read_add(VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z1n6;
wire VMR_L3D3_VMS_L3D3PHI3Z1n6_wr_en;
wire [5:0] VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1_number;
wire [10:0] VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1_read_add;
wire [17:0] VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1;
VMStubs #("Match") VMS_L3D3PHI3Z1n6(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z1n6),
.enable(VMR_L3D3_VMS_L3D3PHI3Z1n6_wr_en),
.number_out(VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1_number),
.read_add(VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1_read_add),
.data_out(VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z2;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2;
VMProjections  VMPROJ_L5L6_L3D3PHI3Z2(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z2),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z2_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2_number),
.read_add(VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D3_VMS_L3D3PHI3Z2n6;
wire VMR_L3D3_VMS_L3D3PHI3Z2n6_wr_en;
wire [5:0] VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2_number;
wire [10:0] VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2_read_add;
wire [17:0] VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2;
VMStubs #("Match") VMS_L3D3PHI3Z2n6(
.data_in(VMR_L3D3_VMS_L3D3PHI3Z2n6),
.enable(VMR_L3D3_VMS_L3D3PHI3Z2n6_wr_en),
.number_out(VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2_number),
.read_add(VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2_read_add),
.data_out(VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z1;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1;
VMProjections  VMPROJ_L5L6_L3D4PHI1Z1(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z1),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z1_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1_number),
.read_add(VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z1n6;
wire VMR_L3D4_VMS_L3D4PHI1Z1n6_wr_en;
wire [5:0] VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1_number;
wire [10:0] VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1_read_add;
wire [17:0] VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1;
VMStubs #("Match") VMS_L3D4PHI1Z1n6(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z1n6),
.enable(VMR_L3D4_VMS_L3D4PHI1Z1n6_wr_en),
.number_out(VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1_number),
.read_add(VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1_read_add),
.data_out(VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z2;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2;
VMProjections  VMPROJ_L5L6_L3D4PHI1Z2(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z2),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z2_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2_number),
.read_add(VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI1Z2n4;
wire VMR_L3D4_VMS_L3D4PHI1Z2n4_wr_en;
wire [5:0] VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2_number;
wire [10:0] VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2_read_add;
wire [17:0] VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2;
VMStubs #("Match") VMS_L3D4PHI1Z2n4(
.data_in(VMR_L3D4_VMS_L3D4PHI1Z2n4),
.enable(VMR_L3D4_VMS_L3D4PHI1Z2n4_wr_en),
.number_out(VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2_number),
.read_add(VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2_read_add),
.data_out(VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z1;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1;
VMProjections  VMPROJ_L5L6_L3D4PHI2Z1(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z1),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z1_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1_number),
.read_add(VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z1n6;
wire VMR_L3D4_VMS_L3D4PHI2Z1n6_wr_en;
wire [5:0] VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1_number;
wire [10:0] VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1_read_add;
wire [17:0] VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1;
VMStubs #("Match") VMS_L3D4PHI2Z1n6(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z1n6),
.enable(VMR_L3D4_VMS_L3D4PHI2Z1n6_wr_en),
.number_out(VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1_number),
.read_add(VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1_read_add),
.data_out(VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z2;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2;
VMProjections  VMPROJ_L5L6_L3D4PHI2Z2(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z2),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z2_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2_number),
.read_add(VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI2Z2n4;
wire VMR_L3D4_VMS_L3D4PHI2Z2n4_wr_en;
wire [5:0] VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2_number;
wire [10:0] VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2_read_add;
wire [17:0] VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2;
VMStubs #("Match") VMS_L3D4PHI2Z2n4(
.data_in(VMR_L3D4_VMS_L3D4PHI2Z2n4),
.enable(VMR_L3D4_VMS_L3D4PHI2Z2n4_wr_en),
.number_out(VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2_number),
.read_add(VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2_read_add),
.data_out(VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z1;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1;
VMProjections  VMPROJ_L5L6_L3D4PHI3Z1(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z1),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z1_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1_number),
.read_add(VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z1n6;
wire VMR_L3D4_VMS_L3D4PHI3Z1n6_wr_en;
wire [5:0] VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1_number;
wire [10:0] VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1_read_add;
wire [17:0] VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1;
VMStubs #("Match") VMS_L3D4PHI3Z1n6(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z1n6),
.enable(VMR_L3D4_VMS_L3D4PHI3Z1n6_wr_en),
.number_out(VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1_number),
.read_add(VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1_read_add),
.data_out(VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z2;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2;
VMProjections  VMPROJ_L5L6_L3D4PHI3Z2(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z2),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z2_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2_number),
.read_add(VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L3D4_VMS_L3D4PHI3Z2n4;
wire VMR_L3D4_VMS_L3D4PHI3Z2n4_wr_en;
wire [5:0] VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2_number;
wire [10:0] VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2_read_add;
wire [17:0] VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2;
VMStubs #("Match") VMS_L3D4PHI3Z2n4(
.data_in(VMR_L3D4_VMS_L3D4PHI3Z2n4),
.enable(VMR_L3D4_VMS_L3D4PHI3Z2n4_wr_en),
.number_out(VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2_number),
.read_add(VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2_read_add),
.data_out(VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z1;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1_read_add;
wire [12:0] VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1;
VMProjections  VMPROJ_L5L6_L4D3PHI1Z1(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z1),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z1_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1_number),
.read_add(VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI1Z1n3;
wire VMR_L4D3_VMS_L4D3PHI1Z1n3_wr_en;
wire [5:0] VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1_number;
wire [10:0] VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1_read_add;
wire [17:0] VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1;
VMStubs #("Match") VMS_L4D3PHI1Z1n3(
.data_in(VMR_L4D3_VMS_L4D3PHI1Z1n3),
.enable(VMR_L4D3_VMS_L4D3PHI1Z1n3_wr_en),
.number_out(VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1_number),
.read_add(VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1_read_add),
.data_out(VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z2;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2_read_add;
wire [12:0] VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2;
VMProjections  VMPROJ_L5L6_L4D3PHI1Z2(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z2),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z2_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2_number),
.read_add(VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI1Z2n4;
wire VMR_L4D3_VMS_L4D3PHI1Z2n4_wr_en;
wire [5:0] VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2_number;
wire [10:0] VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2_read_add;
wire [17:0] VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2;
VMStubs #("Match") VMS_L4D3PHI1Z2n4(
.data_in(VMR_L4D3_VMS_L4D3PHI1Z2n4),
.enable(VMR_L4D3_VMS_L4D3PHI1Z2n4_wr_en),
.number_out(VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2_number),
.read_add(VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2_read_add),
.data_out(VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z1;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1_read_add;
wire [12:0] VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1;
VMProjections  VMPROJ_L5L6_L4D3PHI2Z1(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z1),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z1_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1_number),
.read_add(VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z1n4;
wire VMR_L4D3_VMS_L4D3PHI2Z1n4_wr_en;
wire [5:0] VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1_number;
wire [10:0] VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1_read_add;
wire [17:0] VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1;
VMStubs #("Match") VMS_L4D3PHI2Z1n4(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z1n4),
.enable(VMR_L4D3_VMS_L4D3PHI2Z1n4_wr_en),
.number_out(VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1_number),
.read_add(VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1_read_add),
.data_out(VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z2;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2_read_add;
wire [12:0] VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2;
VMProjections  VMPROJ_L5L6_L4D3PHI2Z2(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z2),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z2_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2_number),
.read_add(VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI2Z2n6;
wire VMR_L4D3_VMS_L4D3PHI2Z2n6_wr_en;
wire [5:0] VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2_number;
wire [10:0] VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2_read_add;
wire [17:0] VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2;
VMStubs #("Match") VMS_L4D3PHI2Z2n6(
.data_in(VMR_L4D3_VMS_L4D3PHI2Z2n6),
.enable(VMR_L4D3_VMS_L4D3PHI2Z2n6_wr_en),
.number_out(VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2_number),
.read_add(VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2_read_add),
.data_out(VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z1;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1_read_add;
wire [12:0] VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1;
VMProjections  VMPROJ_L5L6_L4D3PHI3Z1(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z1),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z1_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1_number),
.read_add(VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z1n4;
wire VMR_L4D3_VMS_L4D3PHI3Z1n4_wr_en;
wire [5:0] VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1_number;
wire [10:0] VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1_read_add;
wire [17:0] VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1;
VMStubs #("Match") VMS_L4D3PHI3Z1n4(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z1n4),
.enable(VMR_L4D3_VMS_L4D3PHI3Z1n4_wr_en),
.number_out(VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1_number),
.read_add(VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1_read_add),
.data_out(VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z2;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2_read_add;
wire [12:0] VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2;
VMProjections  VMPROJ_L5L6_L4D3PHI3Z2(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z2),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z2_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2_number),
.read_add(VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI3Z2n6;
wire VMR_L4D3_VMS_L4D3PHI3Z2n6_wr_en;
wire [5:0] VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2_number;
wire [10:0] VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2_read_add;
wire [17:0] VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2;
VMStubs #("Match") VMS_L4D3PHI3Z2n6(
.data_in(VMR_L4D3_VMS_L4D3PHI3Z2n6),
.enable(VMR_L4D3_VMS_L4D3PHI3Z2n6_wr_en),
.number_out(VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2_number),
.read_add(VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2_read_add),
.data_out(VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z1;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1_read_add;
wire [12:0] VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1;
VMProjections  VMPROJ_L5L6_L4D3PHI4Z1(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z1),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z1_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1_number),
.read_add(VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI4Z1n3;
wire VMR_L4D3_VMS_L4D3PHI4Z1n3_wr_en;
wire [5:0] VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1_number;
wire [10:0] VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1_read_add;
wire [17:0] VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1;
VMStubs #("Match") VMS_L4D3PHI4Z1n3(
.data_in(VMR_L4D3_VMS_L4D3PHI4Z1n3),
.enable(VMR_L4D3_VMS_L4D3PHI4Z1n3_wr_en),
.number_out(VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1_number),
.read_add(VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1_read_add),
.data_out(VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z2;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2_read_add;
wire [12:0] VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2;
VMProjections  VMPROJ_L5L6_L4D3PHI4Z2(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z2),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z2_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2_number),
.read_add(VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D3_VMS_L4D3PHI4Z2n4;
wire VMR_L4D3_VMS_L4D3PHI4Z2n4_wr_en;
wire [5:0] VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2_number;
wire [10:0] VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2_read_add;
wire [17:0] VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2;
VMStubs #("Match") VMS_L4D3PHI4Z2n4(
.data_in(VMR_L4D3_VMS_L4D3PHI4Z2n4),
.enable(VMR_L4D3_VMS_L4D3PHI4Z2n4_wr_en),
.number_out(VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2_number),
.read_add(VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2_read_add),
.data_out(VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z1;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1_read_add;
wire [12:0] VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1;
VMProjections  VMPROJ_L5L6_L4D4PHI1Z1(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z1),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z1_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1_number),
.read_add(VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI1Z1n4;
wire VMR_L4D4_VMS_L4D4PHI1Z1n4_wr_en;
wire [5:0] VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1_number;
wire [10:0] VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1_read_add;
wire [17:0] VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1;
VMStubs #("Match") VMS_L4D4PHI1Z1n4(
.data_in(VMR_L4D4_VMS_L4D4PHI1Z1n4),
.enable(VMR_L4D4_VMS_L4D4PHI1Z1n4_wr_en),
.number_out(VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1_number),
.read_add(VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1_read_add),
.data_out(VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z2;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2_read_add;
wire [12:0] VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2;
VMProjections  VMPROJ_L5L6_L4D4PHI1Z2(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z2),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z2_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2_number),
.read_add(VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI1Z2n4;
wire VMR_L4D4_VMS_L4D4PHI1Z2n4_wr_en;
wire [5:0] VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2_number;
wire [10:0] VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2_read_add;
wire [17:0] VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2;
VMStubs #("Match") VMS_L4D4PHI1Z2n4(
.data_in(VMR_L4D4_VMS_L4D4PHI1Z2n4),
.enable(VMR_L4D4_VMS_L4D4PHI1Z2n4_wr_en),
.number_out(VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2_number),
.read_add(VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2_read_add),
.data_out(VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z1;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1_read_add;
wire [12:0] VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1;
VMProjections  VMPROJ_L5L6_L4D4PHI2Z1(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z1),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z1_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1_number),
.read_add(VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z1n6;
wire VMR_L4D4_VMS_L4D4PHI2Z1n6_wr_en;
wire [5:0] VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1_number;
wire [10:0] VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1_read_add;
wire [17:0] VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1;
VMStubs #("Match") VMS_L4D4PHI2Z1n6(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z1n6),
.enable(VMR_L4D4_VMS_L4D4PHI2Z1n6_wr_en),
.number_out(VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1_number),
.read_add(VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1_read_add),
.data_out(VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z2;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2_read_add;
wire [12:0] VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2;
VMProjections  VMPROJ_L5L6_L4D4PHI2Z2(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z2),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z2_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2_number),
.read_add(VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI2Z2n6;
wire VMR_L4D4_VMS_L4D4PHI2Z2n6_wr_en;
wire [5:0] VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2_number;
wire [10:0] VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2_read_add;
wire [17:0] VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2;
VMStubs #("Match") VMS_L4D4PHI2Z2n6(
.data_in(VMR_L4D4_VMS_L4D4PHI2Z2n6),
.enable(VMR_L4D4_VMS_L4D4PHI2Z2n6_wr_en),
.number_out(VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2_number),
.read_add(VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2_read_add),
.data_out(VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z1;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1_read_add;
wire [12:0] VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1;
VMProjections  VMPROJ_L5L6_L4D4PHI3Z1(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z1),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z1_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1_number),
.read_add(VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z1n6;
wire VMR_L4D4_VMS_L4D4PHI3Z1n6_wr_en;
wire [5:0] VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1_number;
wire [10:0] VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1_read_add;
wire [17:0] VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1;
VMStubs #("Match") VMS_L4D4PHI3Z1n6(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z1n6),
.enable(VMR_L4D4_VMS_L4D4PHI3Z1n6_wr_en),
.number_out(VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1_number),
.read_add(VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1_read_add),
.data_out(VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z2;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2_read_add;
wire [12:0] VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2;
VMProjections  VMPROJ_L5L6_L4D4PHI3Z2(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z2),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z2_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2_number),
.read_add(VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI3Z2n6;
wire VMR_L4D4_VMS_L4D4PHI3Z2n6_wr_en;
wire [5:0] VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2_number;
wire [10:0] VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2_read_add;
wire [17:0] VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2;
VMStubs #("Match") VMS_L4D4PHI3Z2n6(
.data_in(VMR_L4D4_VMS_L4D4PHI3Z2n6),
.enable(VMR_L4D4_VMS_L4D4PHI3Z2n6_wr_en),
.number_out(VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2_number),
.read_add(VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2_read_add),
.data_out(VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z1;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1_read_add;
wire [12:0] VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1;
VMProjections  VMPROJ_L5L6_L4D4PHI4Z1(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z1),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z1_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1_number),
.read_add(VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI4Z1n4;
wire VMR_L4D4_VMS_L4D4PHI4Z1n4_wr_en;
wire [5:0] VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1_number;
wire [10:0] VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1_read_add;
wire [17:0] VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1;
VMStubs #("Match") VMS_L4D4PHI4Z1n4(
.data_in(VMR_L4D4_VMS_L4D4PHI4Z1n4),
.enable(VMR_L4D4_VMS_L4D4PHI4Z1n4_wr_en),
.number_out(VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1_number),
.read_add(VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1_read_add),
.data_out(VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [12:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z2;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2_read_add;
wire [12:0] VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2;
VMProjections  VMPROJ_L5L6_L4D4PHI4Z2(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z2),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z2_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2_number),
.read_add(VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [17:0] VMR_L4D4_VMS_L4D4PHI4Z2n4;
wire VMR_L4D4_VMS_L4D4PHI4Z2n4_wr_en;
wire [5:0] VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2_number;
wire [10:0] VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2_read_add;
wire [17:0] VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2;
VMStubs #("Match") VMS_L4D4PHI4Z2n4(
.data_in(VMR_L4D4_VMS_L4D4PHI4Z2n4),
.enable(VMR_L4D4_VMS_L4D4PHI4Z2n4_wr_en),
.number_out(VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2_number),
.read_add(VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2_read_add),
.data_out(VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D3PHI1Z1_CM_L3L4_L1D3PHI1Z1;
wire ME_L3L4_L1D3PHI1Z1_CM_L3L4_L1D3PHI1Z1_wr_en;
wire [5:0] CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI1Z1(
.data_in(ME_L3L4_L1D3PHI1Z1_CM_L3L4_L1D3PHI1Z1),
.enable(ME_L3L4_L1D3PHI1Z1_CM_L3L4_L1D3PHI1Z1_wr_en),
.number_out(CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3),
.start(start8_0),
.done(done7_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D3PHI1Z2_CM_L3L4_L1D3PHI1Z2;
wire ME_L3L4_L1D3PHI1Z2_CM_L3L4_L1D3PHI1Z2_wr_en;
wire [5:0] CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI1Z2(
.data_in(ME_L3L4_L1D3PHI1Z2_CM_L3L4_L1D3PHI1Z2),
.enable(ME_L3L4_L1D3PHI1Z2_CM_L3L4_L1D3PHI1Z2_wr_en),
.number_out(CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D3PHI2Z1_CM_L3L4_L1D3PHI2Z1;
wire ME_L3L4_L1D3PHI2Z1_CM_L3L4_L1D3PHI2Z1_wr_en;
wire [5:0] CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI2Z1(
.data_in(ME_L3L4_L1D3PHI2Z1_CM_L3L4_L1D3PHI2Z1),
.enable(ME_L3L4_L1D3PHI2Z1_CM_L3L4_L1D3PHI2Z1_wr_en),
.number_out(CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D3PHI2Z2_CM_L3L4_L1D3PHI2Z2;
wire ME_L3L4_L1D3PHI2Z2_CM_L3L4_L1D3PHI2Z2_wr_en;
wire [5:0] CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI2Z2(
.data_in(ME_L3L4_L1D3PHI2Z2_CM_L3L4_L1D3PHI2Z2),
.enable(ME_L3L4_L1D3PHI2Z2_CM_L3L4_L1D3PHI2Z2_wr_en),
.number_out(CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D3PHI3Z1_CM_L3L4_L1D3PHI3Z1;
wire ME_L3L4_L1D3PHI3Z1_CM_L3L4_L1D3PHI3Z1_wr_en;
wire [5:0] CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI3Z1(
.data_in(ME_L3L4_L1D3PHI3Z1_CM_L3L4_L1D3PHI3Z1),
.enable(ME_L3L4_L1D3PHI3Z1_CM_L3L4_L1D3PHI3Z1_wr_en),
.number_out(CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D3PHI3Z2_CM_L3L4_L1D3PHI3Z2;
wire ME_L3L4_L1D3PHI3Z2_CM_L3L4_L1D3PHI3Z2_wr_en;
wire [5:0] CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI3Z2(
.data_in(ME_L3L4_L1D3PHI3Z2_CM_L3L4_L1D3PHI3Z2),
.enable(ME_L3L4_L1D3PHI3Z2_CM_L3L4_L1D3PHI3Z2_wr_en),
.number_out(CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L1D3_L3L4_AP_L3L4_L1D3;
wire PR_L1D3_L3L4_AP_L3L4_L1D3_wr_en;
wire [8:0] AP_L3L4_L1D3_MC_L3L4_L1D3_read_add;
wire [55:0] AP_L3L4_L1D3_MC_L3L4_L1D3;
AllProj #(1'b1) AP_L3L4_L1D3(
.data_in(PR_L1D3_L3L4_AP_L3L4_L1D3),
.enable(PR_L1D3_L3L4_AP_L3L4_L1D3_wr_en),
.read_add(AP_L3L4_L1D3_MC_L3L4_L1D3_read_add),
.data_out(AP_L3L4_L1D3_MC_L3L4_L1D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L1D3_AS_L1D3n3;
wire VMR_L1D3_AS_L1D3n3_wr_en;
wire [10:0] AS_L1D3n3_MC_L3L4_L1D3_read_add;
wire [35:0] AS_L1D3n3_MC_L3L4_L1D3;
AllStubs  AS_L1D3n3(
.data_in(VMR_L1D3_AS_L1D3n3),
.enable(VMR_L1D3_AS_L1D3n3_wr_en),
.read_add_MC(AS_L1D3n3_MC_L3L4_L1D3_read_add),
.data_out_MC(AS_L1D3n3_MC_L3L4_L1D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D4PHI1Z1_CM_L3L4_L1D4PHI1Z1;
wire ME_L3L4_L1D4PHI1Z1_CM_L3L4_L1D4PHI1Z1_wr_en;
wire [5:0] CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI1Z1(
.data_in(ME_L3L4_L1D4PHI1Z1_CM_L3L4_L1D4PHI1Z1),
.enable(ME_L3L4_L1D4PHI1Z1_CM_L3L4_L1D4PHI1Z1_wr_en),
.number_out(CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D4PHI1Z2_CM_L3L4_L1D4PHI1Z2;
wire ME_L3L4_L1D4PHI1Z2_CM_L3L4_L1D4PHI1Z2_wr_en;
wire [5:0] CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI1Z2(
.data_in(ME_L3L4_L1D4PHI1Z2_CM_L3L4_L1D4PHI1Z2),
.enable(ME_L3L4_L1D4PHI1Z2_CM_L3L4_L1D4PHI1Z2_wr_en),
.number_out(CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D4PHI2Z1_CM_L3L4_L1D4PHI2Z1;
wire ME_L3L4_L1D4PHI2Z1_CM_L3L4_L1D4PHI2Z1_wr_en;
wire [5:0] CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI2Z1(
.data_in(ME_L3L4_L1D4PHI2Z1_CM_L3L4_L1D4PHI2Z1),
.enable(ME_L3L4_L1D4PHI2Z1_CM_L3L4_L1D4PHI2Z1_wr_en),
.number_out(CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D4PHI2Z2_CM_L3L4_L1D4PHI2Z2;
wire ME_L3L4_L1D4PHI2Z2_CM_L3L4_L1D4PHI2Z2_wr_en;
wire [5:0] CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI2Z2(
.data_in(ME_L3L4_L1D4PHI2Z2_CM_L3L4_L1D4PHI2Z2),
.enable(ME_L3L4_L1D4PHI2Z2_CM_L3L4_L1D4PHI2Z2_wr_en),
.number_out(CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D4PHI3Z1_CM_L3L4_L1D4PHI3Z1;
wire ME_L3L4_L1D4PHI3Z1_CM_L3L4_L1D4PHI3Z1_wr_en;
wire [5:0] CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI3Z1(
.data_in(ME_L3L4_L1D4PHI3Z1_CM_L3L4_L1D4PHI3Z1),
.enable(ME_L3L4_L1D4PHI3Z1_CM_L3L4_L1D4PHI3Z1_wr_en),
.number_out(CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L1D4PHI3Z2_CM_L3L4_L1D4PHI3Z2;
wire ME_L3L4_L1D4PHI3Z2_CM_L3L4_L1D4PHI3Z2_wr_en;
wire [5:0] CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI3Z2(
.data_in(ME_L3L4_L1D4PHI3Z2_CM_L3L4_L1D4PHI3Z2),
.enable(ME_L3L4_L1D4PHI3Z2_CM_L3L4_L1D4PHI3Z2_wr_en),
.number_out(CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L1D4_L3L4_AP_L3L4_L1D4;
wire PR_L1D4_L3L4_AP_L3L4_L1D4_wr_en;
wire [8:0] AP_L3L4_L1D4_MC_L3L4_L1D4_read_add;
wire [55:0] AP_L3L4_L1D4_MC_L3L4_L1D4;
AllProj #(1'b1) AP_L3L4_L1D4(
.data_in(PR_L1D4_L3L4_AP_L3L4_L1D4),
.enable(PR_L1D4_L3L4_AP_L3L4_L1D4_wr_en),
.read_add(AP_L3L4_L1D4_MC_L3L4_L1D4_read_add),
.data_out(AP_L3L4_L1D4_MC_L3L4_L1D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L1D4_AS_L1D4n2;
wire VMR_L1D4_AS_L1D4n2_wr_en;
wire [10:0] AS_L1D4n2_MC_L3L4_L1D4_read_add;
wire [35:0] AS_L1D4n2_MC_L3L4_L1D4;
AllStubs  AS_L1D4n2(
.data_in(VMR_L1D4_AS_L1D4n2),
.enable(VMR_L1D4_AS_L1D4n2_wr_en),
.read_add_MC(AS_L1D4n2_MC_L3L4_L1D4_read_add),
.data_out_MC(AS_L1D4n2_MC_L3L4_L1D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D3PHI1Z1_CM_L3L4_L2D3PHI1Z1;
wire ME_L3L4_L2D3PHI1Z1_CM_L3L4_L2D3PHI1Z1_wr_en;
wire [5:0] CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI1Z1(
.data_in(ME_L3L4_L2D3PHI1Z1_CM_L3L4_L2D3PHI1Z1),
.enable(ME_L3L4_L2D3PHI1Z1_CM_L3L4_L2D3PHI1Z1_wr_en),
.number_out(CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D3PHI1Z2_CM_L3L4_L2D3PHI1Z2;
wire ME_L3L4_L2D3PHI1Z2_CM_L3L4_L2D3PHI1Z2_wr_en;
wire [5:0] CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI1Z2(
.data_in(ME_L3L4_L2D3PHI1Z2_CM_L3L4_L2D3PHI1Z2),
.enable(ME_L3L4_L2D3PHI1Z2_CM_L3L4_L2D3PHI1Z2_wr_en),
.number_out(CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D3PHI2Z1_CM_L3L4_L2D3PHI2Z1;
wire ME_L3L4_L2D3PHI2Z1_CM_L3L4_L2D3PHI2Z1_wr_en;
wire [5:0] CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI2Z1(
.data_in(ME_L3L4_L2D3PHI2Z1_CM_L3L4_L2D3PHI2Z1),
.enable(ME_L3L4_L2D3PHI2Z1_CM_L3L4_L2D3PHI2Z1_wr_en),
.number_out(CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D3PHI2Z2_CM_L3L4_L2D3PHI2Z2;
wire ME_L3L4_L2D3PHI2Z2_CM_L3L4_L2D3PHI2Z2_wr_en;
wire [5:0] CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI2Z2(
.data_in(ME_L3L4_L2D3PHI2Z2_CM_L3L4_L2D3PHI2Z2),
.enable(ME_L3L4_L2D3PHI2Z2_CM_L3L4_L2D3PHI2Z2_wr_en),
.number_out(CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D3PHI3Z1_CM_L3L4_L2D3PHI3Z1;
wire ME_L3L4_L2D3PHI3Z1_CM_L3L4_L2D3PHI3Z1_wr_en;
wire [5:0] CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI3Z1(
.data_in(ME_L3L4_L2D3PHI3Z1_CM_L3L4_L2D3PHI3Z1),
.enable(ME_L3L4_L2D3PHI3Z1_CM_L3L4_L2D3PHI3Z1_wr_en),
.number_out(CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D3PHI3Z2_CM_L3L4_L2D3PHI3Z2;
wire ME_L3L4_L2D3PHI3Z2_CM_L3L4_L2D3PHI3Z2_wr_en;
wire [5:0] CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI3Z2(
.data_in(ME_L3L4_L2D3PHI3Z2_CM_L3L4_L2D3PHI3Z2),
.enable(ME_L3L4_L2D3PHI3Z2_CM_L3L4_L2D3PHI3Z2_wr_en),
.number_out(CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D3PHI4Z1_CM_L3L4_L2D3PHI4Z1;
wire ME_L3L4_L2D3PHI4Z1_CM_L3L4_L2D3PHI4Z1_wr_en;
wire [5:0] CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI4Z1(
.data_in(ME_L3L4_L2D3PHI4Z1_CM_L3L4_L2D3PHI4Z1),
.enable(ME_L3L4_L2D3PHI4Z1_CM_L3L4_L2D3PHI4Z1_wr_en),
.number_out(CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D3PHI4Z2_CM_L3L4_L2D3PHI4Z2;
wire ME_L3L4_L2D3PHI4Z2_CM_L3L4_L2D3PHI4Z2_wr_en;
wire [5:0] CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI4Z2(
.data_in(ME_L3L4_L2D3PHI4Z2_CM_L3L4_L2D3PHI4Z2),
.enable(ME_L3L4_L2D3PHI4Z2_CM_L3L4_L2D3PHI4Z2_wr_en),
.number_out(CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L2D3_L3L4_AP_L3L4_L2D3;
wire PR_L2D3_L3L4_AP_L3L4_L2D3_wr_en;
wire [8:0] AP_L3L4_L2D3_MC_L3L4_L2D3_read_add;
wire [55:0] AP_L3L4_L2D3_MC_L3L4_L2D3;
AllProj #(1'b1) AP_L3L4_L2D3(
.data_in(PR_L2D3_L3L4_AP_L3L4_L2D3),
.enable(PR_L2D3_L3L4_AP_L3L4_L2D3_wr_en),
.read_add(AP_L3L4_L2D3_MC_L3L4_L2D3_read_add),
.data_out(AP_L3L4_L2D3_MC_L3L4_L2D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L2D3_AS_L2D3n2;
wire VMR_L2D3_AS_L2D3n2_wr_en;
wire [10:0] AS_L2D3n2_MC_L3L4_L2D3_read_add;
wire [35:0] AS_L2D3n2_MC_L3L4_L2D3;
AllStubs  AS_L2D3n2(
.data_in(VMR_L2D3_AS_L2D3n2),
.enable(VMR_L2D3_AS_L2D3n2_wr_en),
.read_add_MC(AS_L2D3n2_MC_L3L4_L2D3_read_add),
.data_out_MC(AS_L2D3n2_MC_L3L4_L2D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D4PHI1Z1_CM_L3L4_L2D4PHI1Z1;
wire ME_L3L4_L2D4PHI1Z1_CM_L3L4_L2D4PHI1Z1_wr_en;
wire [5:0] CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI1Z1(
.data_in(ME_L3L4_L2D4PHI1Z1_CM_L3L4_L2D4PHI1Z1),
.enable(ME_L3L4_L2D4PHI1Z1_CM_L3L4_L2D4PHI1Z1_wr_en),
.number_out(CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D4PHI1Z2_CM_L3L4_L2D4PHI1Z2;
wire ME_L3L4_L2D4PHI1Z2_CM_L3L4_L2D4PHI1Z2_wr_en;
wire [5:0] CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI1Z2(
.data_in(ME_L3L4_L2D4PHI1Z2_CM_L3L4_L2D4PHI1Z2),
.enable(ME_L3L4_L2D4PHI1Z2_CM_L3L4_L2D4PHI1Z2_wr_en),
.number_out(CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D4PHI2Z1_CM_L3L4_L2D4PHI2Z1;
wire ME_L3L4_L2D4PHI2Z1_CM_L3L4_L2D4PHI2Z1_wr_en;
wire [5:0] CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI2Z1(
.data_in(ME_L3L4_L2D4PHI2Z1_CM_L3L4_L2D4PHI2Z1),
.enable(ME_L3L4_L2D4PHI2Z1_CM_L3L4_L2D4PHI2Z1_wr_en),
.number_out(CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D4PHI2Z2_CM_L3L4_L2D4PHI2Z2;
wire ME_L3L4_L2D4PHI2Z2_CM_L3L4_L2D4PHI2Z2_wr_en;
wire [5:0] CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI2Z2(
.data_in(ME_L3L4_L2D4PHI2Z2_CM_L3L4_L2D4PHI2Z2),
.enable(ME_L3L4_L2D4PHI2Z2_CM_L3L4_L2D4PHI2Z2_wr_en),
.number_out(CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D4PHI3Z1_CM_L3L4_L2D4PHI3Z1;
wire ME_L3L4_L2D4PHI3Z1_CM_L3L4_L2D4PHI3Z1_wr_en;
wire [5:0] CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI3Z1(
.data_in(ME_L3L4_L2D4PHI3Z1_CM_L3L4_L2D4PHI3Z1),
.enable(ME_L3L4_L2D4PHI3Z1_CM_L3L4_L2D4PHI3Z1_wr_en),
.number_out(CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D4PHI3Z2_CM_L3L4_L2D4PHI3Z2;
wire ME_L3L4_L2D4PHI3Z2_CM_L3L4_L2D4PHI3Z2_wr_en;
wire [5:0] CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI3Z2(
.data_in(ME_L3L4_L2D4PHI3Z2_CM_L3L4_L2D4PHI3Z2),
.enable(ME_L3L4_L2D4PHI3Z2_CM_L3L4_L2D4PHI3Z2_wr_en),
.number_out(CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D4PHI4Z1_CM_L3L4_L2D4PHI4Z1;
wire ME_L3L4_L2D4PHI4Z1_CM_L3L4_L2D4PHI4Z1_wr_en;
wire [5:0] CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI4Z1(
.data_in(ME_L3L4_L2D4PHI4Z1_CM_L3L4_L2D4PHI4Z1),
.enable(ME_L3L4_L2D4PHI4Z1_CM_L3L4_L2D4PHI4Z1_wr_en),
.number_out(CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L2D4PHI4Z2_CM_L3L4_L2D4PHI4Z2;
wire ME_L3L4_L2D4PHI4Z2_CM_L3L4_L2D4PHI4Z2_wr_en;
wire [5:0] CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI4Z2(
.data_in(ME_L3L4_L2D4PHI4Z2_CM_L3L4_L2D4PHI4Z2),
.enable(ME_L3L4_L2D4PHI4Z2_CM_L3L4_L2D4PHI4Z2_wr_en),
.number_out(CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L2D4_L3L4_AP_L3L4_L2D4;
wire PR_L2D4_L3L4_AP_L3L4_L2D4_wr_en;
wire [8:0] AP_L3L4_L2D4_MC_L3L4_L2D4_read_add;
wire [55:0] AP_L3L4_L2D4_MC_L3L4_L2D4;
AllProj #(1'b1) AP_L3L4_L2D4(
.data_in(PR_L2D4_L3L4_AP_L3L4_L2D4),
.enable(PR_L2D4_L3L4_AP_L3L4_L2D4_wr_en),
.read_add(AP_L3L4_L2D4_MC_L3L4_L2D4_read_add),
.data_out(AP_L3L4_L2D4_MC_L3L4_L2D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L2D4_AS_L2D4n3;
wire VMR_L2D4_AS_L2D4n3_wr_en;
wire [10:0] AS_L2D4n3_MC_L3L4_L2D4_read_add;
wire [35:0] AS_L2D4n3_MC_L3L4_L2D4;
AllStubs  AS_L2D4n3(
.data_in(VMR_L2D4_AS_L2D4n3),
.enable(VMR_L2D4_AS_L2D4n3_wr_en),
.read_add_MC(AS_L2D4n3_MC_L3L4_L2D4_read_add),
.data_out_MC(AS_L2D4n3_MC_L3L4_L2D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D3PHI1Z1_CM_L3L4_L5D3PHI1Z1;
wire ME_L3L4_L5D3PHI1Z1_CM_L3L4_L5D3PHI1Z1_wr_en;
wire [5:0] CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI1Z1(
.data_in(ME_L3L4_L5D3PHI1Z1_CM_L3L4_L5D3PHI1Z1),
.enable(ME_L3L4_L5D3PHI1Z1_CM_L3L4_L5D3PHI1Z1_wr_en),
.number_out(CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D3PHI1Z2_CM_L3L4_L5D3PHI1Z2;
wire ME_L3L4_L5D3PHI1Z2_CM_L3L4_L5D3PHI1Z2_wr_en;
wire [5:0] CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI1Z2(
.data_in(ME_L3L4_L5D3PHI1Z2_CM_L3L4_L5D3PHI1Z2),
.enable(ME_L3L4_L5D3PHI1Z2_CM_L3L4_L5D3PHI1Z2_wr_en),
.number_out(CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D3PHI2Z1_CM_L3L4_L5D3PHI2Z1;
wire ME_L3L4_L5D3PHI2Z1_CM_L3L4_L5D3PHI2Z1_wr_en;
wire [5:0] CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI2Z1(
.data_in(ME_L3L4_L5D3PHI2Z1_CM_L3L4_L5D3PHI2Z1),
.enable(ME_L3L4_L5D3PHI2Z1_CM_L3L4_L5D3PHI2Z1_wr_en),
.number_out(CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D3PHI2Z2_CM_L3L4_L5D3PHI2Z2;
wire ME_L3L4_L5D3PHI2Z2_CM_L3L4_L5D3PHI2Z2_wr_en;
wire [5:0] CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI2Z2(
.data_in(ME_L3L4_L5D3PHI2Z2_CM_L3L4_L5D3PHI2Z2),
.enable(ME_L3L4_L5D3PHI2Z2_CM_L3L4_L5D3PHI2Z2_wr_en),
.number_out(CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D3PHI3Z1_CM_L3L4_L5D3PHI3Z1;
wire ME_L3L4_L5D3PHI3Z1_CM_L3L4_L5D3PHI3Z1_wr_en;
wire [5:0] CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI3Z1(
.data_in(ME_L3L4_L5D3PHI3Z1_CM_L3L4_L5D3PHI3Z1),
.enable(ME_L3L4_L5D3PHI3Z1_CM_L3L4_L5D3PHI3Z1_wr_en),
.number_out(CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D3PHI3Z2_CM_L3L4_L5D3PHI3Z2;
wire ME_L3L4_L5D3PHI3Z2_CM_L3L4_L5D3PHI3Z2_wr_en;
wire [5:0] CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI3Z2(
.data_in(ME_L3L4_L5D3PHI3Z2_CM_L3L4_L5D3PHI3Z2),
.enable(ME_L3L4_L5D3PHI3Z2_CM_L3L4_L5D3PHI3Z2_wr_en),
.number_out(CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L5D3_L3L4_AP_L3L4_L5D3;
wire PR_L5D3_L3L4_AP_L3L4_L5D3_wr_en;
wire [8:0] AP_L3L4_L5D3_MC_L3L4_L5D3_read_add;
wire [55:0] AP_L3L4_L5D3_MC_L3L4_L5D3;
AllProj #(1'b0) AP_L3L4_L5D3(
.data_in(PR_L5D3_L3L4_AP_L3L4_L5D3),
.enable(PR_L5D3_L3L4_AP_L3L4_L5D3_wr_en),
.read_add(AP_L3L4_L5D3_MC_L3L4_L5D3_read_add),
.data_out(AP_L3L4_L5D3_MC_L3L4_L5D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L5D3_AS_L5D3n3;
wire VMR_L5D3_AS_L5D3n3_wr_en;
wire [10:0] AS_L5D3n3_MC_L3L4_L5D3_read_add;
wire [35:0] AS_L5D3n3_MC_L3L4_L5D3;
AllStubs  AS_L5D3n3(
.data_in(VMR_L5D3_AS_L5D3n3),
.enable(VMR_L5D3_AS_L5D3n3_wr_en),
.read_add_MC(AS_L5D3n3_MC_L3L4_L5D3_read_add),
.data_out_MC(AS_L5D3n3_MC_L3L4_L5D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D4PHI1Z1_CM_L3L4_L5D4PHI1Z1;
wire ME_L3L4_L5D4PHI1Z1_CM_L3L4_L5D4PHI1Z1_wr_en;
wire [5:0] CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI1Z1(
.data_in(ME_L3L4_L5D4PHI1Z1_CM_L3L4_L5D4PHI1Z1),
.enable(ME_L3L4_L5D4PHI1Z1_CM_L3L4_L5D4PHI1Z1_wr_en),
.number_out(CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D4PHI1Z2_CM_L3L4_L5D4PHI1Z2;
wire ME_L3L4_L5D4PHI1Z2_CM_L3L4_L5D4PHI1Z2_wr_en;
wire [5:0] CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI1Z2(
.data_in(ME_L3L4_L5D4PHI1Z2_CM_L3L4_L5D4PHI1Z2),
.enable(ME_L3L4_L5D4PHI1Z2_CM_L3L4_L5D4PHI1Z2_wr_en),
.number_out(CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D4PHI2Z1_CM_L3L4_L5D4PHI2Z1;
wire ME_L3L4_L5D4PHI2Z1_CM_L3L4_L5D4PHI2Z1_wr_en;
wire [5:0] CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI2Z1(
.data_in(ME_L3L4_L5D4PHI2Z1_CM_L3L4_L5D4PHI2Z1),
.enable(ME_L3L4_L5D4PHI2Z1_CM_L3L4_L5D4PHI2Z1_wr_en),
.number_out(CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D4PHI2Z2_CM_L3L4_L5D4PHI2Z2;
wire ME_L3L4_L5D4PHI2Z2_CM_L3L4_L5D4PHI2Z2_wr_en;
wire [5:0] CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI2Z2(
.data_in(ME_L3L4_L5D4PHI2Z2_CM_L3L4_L5D4PHI2Z2),
.enable(ME_L3L4_L5D4PHI2Z2_CM_L3L4_L5D4PHI2Z2_wr_en),
.number_out(CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D4PHI3Z1_CM_L3L4_L5D4PHI3Z1;
wire ME_L3L4_L5D4PHI3Z1_CM_L3L4_L5D4PHI3Z1_wr_en;
wire [5:0] CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI3Z1(
.data_in(ME_L3L4_L5D4PHI3Z1_CM_L3L4_L5D4PHI3Z1),
.enable(ME_L3L4_L5D4PHI3Z1_CM_L3L4_L5D4PHI3Z1_wr_en),
.number_out(CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L5D4PHI3Z2_CM_L3L4_L5D4PHI3Z2;
wire ME_L3L4_L5D4PHI3Z2_CM_L3L4_L5D4PHI3Z2_wr_en;
wire [5:0] CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI3Z2(
.data_in(ME_L3L4_L5D4PHI3Z2_CM_L3L4_L5D4PHI3Z2),
.enable(ME_L3L4_L5D4PHI3Z2_CM_L3L4_L5D4PHI3Z2_wr_en),
.number_out(CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L5D4_L3L4_AP_L3L4_L5D4;
wire PR_L5D4_L3L4_AP_L3L4_L5D4_wr_en;
wire [8:0] AP_L3L4_L5D4_MC_L3L4_L5D4_read_add;
wire [55:0] AP_L3L4_L5D4_MC_L3L4_L5D4;
AllProj #(1'b0) AP_L3L4_L5D4(
.data_in(PR_L5D4_L3L4_AP_L3L4_L5D4),
.enable(PR_L5D4_L3L4_AP_L3L4_L5D4_wr_en),
.read_add(AP_L3L4_L5D4_MC_L3L4_L5D4_read_add),
.data_out(AP_L3L4_L5D4_MC_L3L4_L5D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L5D4_AS_L5D4n2;
wire VMR_L5D4_AS_L5D4n2_wr_en;
wire [10:0] AS_L5D4n2_MC_L3L4_L5D4_read_add;
wire [35:0] AS_L5D4n2_MC_L3L4_L5D4;
AllStubs  AS_L5D4n2(
.data_in(VMR_L5D4_AS_L5D4n2),
.enable(VMR_L5D4_AS_L5D4n2_wr_en),
.read_add_MC(AS_L5D4n2_MC_L3L4_L5D4_read_add),
.data_out_MC(AS_L5D4n2_MC_L3L4_L5D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D3PHI1Z1_CM_L3L4_L6D3PHI1Z1;
wire ME_L3L4_L6D3PHI1Z1_CM_L3L4_L6D3PHI1Z1_wr_en;
wire [5:0] CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI1Z1(
.data_in(ME_L3L4_L6D3PHI1Z1_CM_L3L4_L6D3PHI1Z1),
.enable(ME_L3L4_L6D3PHI1Z1_CM_L3L4_L6D3PHI1Z1_wr_en),
.number_out(CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D3PHI1Z2_CM_L3L4_L6D3PHI1Z2;
wire ME_L3L4_L6D3PHI1Z2_CM_L3L4_L6D3PHI1Z2_wr_en;
wire [5:0] CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI1Z2(
.data_in(ME_L3L4_L6D3PHI1Z2_CM_L3L4_L6D3PHI1Z2),
.enable(ME_L3L4_L6D3PHI1Z2_CM_L3L4_L6D3PHI1Z2_wr_en),
.number_out(CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D3PHI2Z1_CM_L3L4_L6D3PHI2Z1;
wire ME_L3L4_L6D3PHI2Z1_CM_L3L4_L6D3PHI2Z1_wr_en;
wire [5:0] CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI2Z1(
.data_in(ME_L3L4_L6D3PHI2Z1_CM_L3L4_L6D3PHI2Z1),
.enable(ME_L3L4_L6D3PHI2Z1_CM_L3L4_L6D3PHI2Z1_wr_en),
.number_out(CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D3PHI2Z2_CM_L3L4_L6D3PHI2Z2;
wire ME_L3L4_L6D3PHI2Z2_CM_L3L4_L6D3PHI2Z2_wr_en;
wire [5:0] CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI2Z2(
.data_in(ME_L3L4_L6D3PHI2Z2_CM_L3L4_L6D3PHI2Z2),
.enable(ME_L3L4_L6D3PHI2Z2_CM_L3L4_L6D3PHI2Z2_wr_en),
.number_out(CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D3PHI3Z1_CM_L3L4_L6D3PHI3Z1;
wire ME_L3L4_L6D3PHI3Z1_CM_L3L4_L6D3PHI3Z1_wr_en;
wire [5:0] CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI3Z1(
.data_in(ME_L3L4_L6D3PHI3Z1_CM_L3L4_L6D3PHI3Z1),
.enable(ME_L3L4_L6D3PHI3Z1_CM_L3L4_L6D3PHI3Z1_wr_en),
.number_out(CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D3PHI3Z2_CM_L3L4_L6D3PHI3Z2;
wire ME_L3L4_L6D3PHI3Z2_CM_L3L4_L6D3PHI3Z2_wr_en;
wire [5:0] CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI3Z2(
.data_in(ME_L3L4_L6D3PHI3Z2_CM_L3L4_L6D3PHI3Z2),
.enable(ME_L3L4_L6D3PHI3Z2_CM_L3L4_L6D3PHI3Z2_wr_en),
.number_out(CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D3PHI4Z1_CM_L3L4_L6D3PHI4Z1;
wire ME_L3L4_L6D3PHI4Z1_CM_L3L4_L6D3PHI4Z1_wr_en;
wire [5:0] CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI4Z1(
.data_in(ME_L3L4_L6D3PHI4Z1_CM_L3L4_L6D3PHI4Z1),
.enable(ME_L3L4_L6D3PHI4Z1_CM_L3L4_L6D3PHI4Z1_wr_en),
.number_out(CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D3PHI4Z2_CM_L3L4_L6D3PHI4Z2;
wire ME_L3L4_L6D3PHI4Z2_CM_L3L4_L6D3PHI4Z2_wr_en;
wire [5:0] CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI4Z2(
.data_in(ME_L3L4_L6D3PHI4Z2_CM_L3L4_L6D3PHI4Z2),
.enable(ME_L3L4_L6D3PHI4Z2_CM_L3L4_L6D3PHI4Z2_wr_en),
.number_out(CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L6D3_L3L4_AP_L3L4_L6D3;
wire PR_L6D3_L3L4_AP_L3L4_L6D3_wr_en;
wire [8:0] AP_L3L4_L6D3_MC_L3L4_L6D3_read_add;
wire [55:0] AP_L3L4_L6D3_MC_L3L4_L6D3;
AllProj #(1'b0) AP_L3L4_L6D3(
.data_in(PR_L6D3_L3L4_AP_L3L4_L6D3),
.enable(PR_L6D3_L3L4_AP_L3L4_L6D3_wr_en),
.read_add(AP_L3L4_L6D3_MC_L3L4_L6D3_read_add),
.data_out(AP_L3L4_L6D3_MC_L3L4_L6D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L6D3_AS_L6D3n2;
wire VMR_L6D3_AS_L6D3n2_wr_en;
wire [10:0] AS_L6D3n2_MC_L3L4_L6D3_read_add;
wire [35:0] AS_L6D3n2_MC_L3L4_L6D3;
AllStubs  AS_L6D3n2(
.data_in(VMR_L6D3_AS_L6D3n2),
.enable(VMR_L6D3_AS_L6D3n2_wr_en),
.read_add_MC(AS_L6D3n2_MC_L3L4_L6D3_read_add),
.data_out_MC(AS_L6D3n2_MC_L3L4_L6D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D4PHI1Z1_CM_L3L4_L6D4PHI1Z1;
wire ME_L3L4_L6D4PHI1Z1_CM_L3L4_L6D4PHI1Z1_wr_en;
wire [5:0] CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI1Z1(
.data_in(ME_L3L4_L6D4PHI1Z1_CM_L3L4_L6D4PHI1Z1),
.enable(ME_L3L4_L6D4PHI1Z1_CM_L3L4_L6D4PHI1Z1_wr_en),
.number_out(CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D4PHI1Z2_CM_L3L4_L6D4PHI1Z2;
wire ME_L3L4_L6D4PHI1Z2_CM_L3L4_L6D4PHI1Z2_wr_en;
wire [5:0] CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI1Z2(
.data_in(ME_L3L4_L6D4PHI1Z2_CM_L3L4_L6D4PHI1Z2),
.enable(ME_L3L4_L6D4PHI1Z2_CM_L3L4_L6D4PHI1Z2_wr_en),
.number_out(CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D4PHI2Z1_CM_L3L4_L6D4PHI2Z1;
wire ME_L3L4_L6D4PHI2Z1_CM_L3L4_L6D4PHI2Z1_wr_en;
wire [5:0] CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI2Z1(
.data_in(ME_L3L4_L6D4PHI2Z1_CM_L3L4_L6D4PHI2Z1),
.enable(ME_L3L4_L6D4PHI2Z1_CM_L3L4_L6D4PHI2Z1_wr_en),
.number_out(CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D4PHI2Z2_CM_L3L4_L6D4PHI2Z2;
wire ME_L3L4_L6D4PHI2Z2_CM_L3L4_L6D4PHI2Z2_wr_en;
wire [5:0] CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI2Z2(
.data_in(ME_L3L4_L6D4PHI2Z2_CM_L3L4_L6D4PHI2Z2),
.enable(ME_L3L4_L6D4PHI2Z2_CM_L3L4_L6D4PHI2Z2_wr_en),
.number_out(CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D4PHI3Z1_CM_L3L4_L6D4PHI3Z1;
wire ME_L3L4_L6D4PHI3Z1_CM_L3L4_L6D4PHI3Z1_wr_en;
wire [5:0] CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI3Z1(
.data_in(ME_L3L4_L6D4PHI3Z1_CM_L3L4_L6D4PHI3Z1),
.enable(ME_L3L4_L6D4PHI3Z1_CM_L3L4_L6D4PHI3Z1_wr_en),
.number_out(CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D4PHI3Z2_CM_L3L4_L6D4PHI3Z2;
wire ME_L3L4_L6D4PHI3Z2_CM_L3L4_L6D4PHI3Z2_wr_en;
wire [5:0] CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI3Z2(
.data_in(ME_L3L4_L6D4PHI3Z2_CM_L3L4_L6D4PHI3Z2),
.enable(ME_L3L4_L6D4PHI3Z2_CM_L3L4_L6D4PHI3Z2_wr_en),
.number_out(CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D4PHI4Z1_CM_L3L4_L6D4PHI4Z1;
wire ME_L3L4_L6D4PHI4Z1_CM_L3L4_L6D4PHI4Z1_wr_en;
wire [5:0] CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI4Z1(
.data_in(ME_L3L4_L6D4PHI4Z1_CM_L3L4_L6D4PHI4Z1),
.enable(ME_L3L4_L6D4PHI4Z1_CM_L3L4_L6D4PHI4Z1_wr_en),
.number_out(CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L3L4_L6D4PHI4Z2_CM_L3L4_L6D4PHI4Z2;
wire ME_L3L4_L6D4PHI4Z2_CM_L3L4_L6D4PHI4Z2_wr_en;
wire [5:0] CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI4Z2(
.data_in(ME_L3L4_L6D4PHI4Z2_CM_L3L4_L6D4PHI4Z2),
.enable(ME_L3L4_L6D4PHI4Z2_CM_L3L4_L6D4PHI4Z2_wr_en),
.number_out(CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L6D4_L3L4_AP_L3L4_L6D4;
wire PR_L6D4_L3L4_AP_L3L4_L6D4_wr_en;
wire [8:0] AP_L3L4_L6D4_MC_L3L4_L6D4_read_add;
wire [55:0] AP_L3L4_L6D4_MC_L3L4_L6D4;
AllProj #(1'b0) AP_L3L4_L6D4(
.data_in(PR_L6D4_L3L4_AP_L3L4_L6D4),
.enable(PR_L6D4_L3L4_AP_L3L4_L6D4_wr_en),
.read_add(AP_L3L4_L6D4_MC_L3L4_L6D4_read_add),
.data_out(AP_L3L4_L6D4_MC_L3L4_L6D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L6D4_AS_L6D4n3;
wire VMR_L6D4_AS_L6D4n3_wr_en;
wire [10:0] AS_L6D4n3_MC_L3L4_L6D4_read_add;
wire [35:0] AS_L6D4n3_MC_L3L4_L6D4;
AllStubs  AS_L6D4n3(
.data_in(VMR_L6D4_AS_L6D4n3),
.enable(VMR_L6D4_AS_L6D4n3_wr_en),
.read_add_MC(AS_L6D4n3_MC_L3L4_L6D4_read_add),
.data_out_MC(AS_L6D4n3_MC_L3L4_L6D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D3PHI1Z1_CM_L5L6_L1D3PHI1Z1;
wire ME_L5L6_L1D3PHI1Z1_CM_L5L6_L1D3PHI1Z1_wr_en;
wire [5:0] CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI1Z1(
.data_in(ME_L5L6_L1D3PHI1Z1_CM_L5L6_L1D3PHI1Z1),
.enable(ME_L5L6_L1D3PHI1Z1_CM_L5L6_L1D3PHI1Z1_wr_en),
.number_out(CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D3PHI1Z2_CM_L5L6_L1D3PHI1Z2;
wire ME_L5L6_L1D3PHI1Z2_CM_L5L6_L1D3PHI1Z2_wr_en;
wire [5:0] CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI1Z2(
.data_in(ME_L5L6_L1D3PHI1Z2_CM_L5L6_L1D3PHI1Z2),
.enable(ME_L5L6_L1D3PHI1Z2_CM_L5L6_L1D3PHI1Z2_wr_en),
.number_out(CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D3PHI2Z1_CM_L5L6_L1D3PHI2Z1;
wire ME_L5L6_L1D3PHI2Z1_CM_L5L6_L1D3PHI2Z1_wr_en;
wire [5:0] CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI2Z1(
.data_in(ME_L5L6_L1D3PHI2Z1_CM_L5L6_L1D3PHI2Z1),
.enable(ME_L5L6_L1D3PHI2Z1_CM_L5L6_L1D3PHI2Z1_wr_en),
.number_out(CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D3PHI2Z2_CM_L5L6_L1D3PHI2Z2;
wire ME_L5L6_L1D3PHI2Z2_CM_L5L6_L1D3PHI2Z2_wr_en;
wire [5:0] CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI2Z2(
.data_in(ME_L5L6_L1D3PHI2Z2_CM_L5L6_L1D3PHI2Z2),
.enable(ME_L5L6_L1D3PHI2Z2_CM_L5L6_L1D3PHI2Z2_wr_en),
.number_out(CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D3PHI3Z1_CM_L5L6_L1D3PHI3Z1;
wire ME_L5L6_L1D3PHI3Z1_CM_L5L6_L1D3PHI3Z1_wr_en;
wire [5:0] CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI3Z1(
.data_in(ME_L5L6_L1D3PHI3Z1_CM_L5L6_L1D3PHI3Z1),
.enable(ME_L5L6_L1D3PHI3Z1_CM_L5L6_L1D3PHI3Z1_wr_en),
.number_out(CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D3PHI3Z2_CM_L5L6_L1D3PHI3Z2;
wire ME_L5L6_L1D3PHI3Z2_CM_L5L6_L1D3PHI3Z2_wr_en;
wire [5:0] CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI3Z2(
.data_in(ME_L5L6_L1D3PHI3Z2_CM_L5L6_L1D3PHI3Z2),
.enable(ME_L5L6_L1D3PHI3Z2_CM_L5L6_L1D3PHI3Z2_wr_en),
.number_out(CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L1D3_L5L6_AP_L5L6_L1D3;
wire PR_L1D3_L5L6_AP_L5L6_L1D3_wr_en;
wire [8:0] AP_L5L6_L1D3_MC_L5L6_L1D3_read_add;
wire [55:0] AP_L5L6_L1D3_MC_L5L6_L1D3;
AllProj #(1'b1) AP_L5L6_L1D3(
.data_in(PR_L1D3_L5L6_AP_L5L6_L1D3),
.enable(PR_L1D3_L5L6_AP_L5L6_L1D3_wr_en),
.read_add(AP_L5L6_L1D3_MC_L5L6_L1D3_read_add),
.data_out(AP_L5L6_L1D3_MC_L5L6_L1D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L1D3_AS_L1D3n4;
wire VMR_L1D3_AS_L1D3n4_wr_en;
wire [10:0] AS_L1D3n4_MC_L5L6_L1D3_read_add;
wire [35:0] AS_L1D3n4_MC_L5L6_L1D3;
AllStubs  AS_L1D3n4(
.data_in(VMR_L1D3_AS_L1D3n4),
.enable(VMR_L1D3_AS_L1D3n4_wr_en),
.read_add_MC(AS_L1D3n4_MC_L5L6_L1D3_read_add),
.data_out_MC(AS_L1D3n4_MC_L5L6_L1D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D4PHI1Z1_CM_L5L6_L1D4PHI1Z1;
wire ME_L5L6_L1D4PHI1Z1_CM_L5L6_L1D4PHI1Z1_wr_en;
wire [5:0] CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI1Z1(
.data_in(ME_L5L6_L1D4PHI1Z1_CM_L5L6_L1D4PHI1Z1),
.enable(ME_L5L6_L1D4PHI1Z1_CM_L5L6_L1D4PHI1Z1_wr_en),
.number_out(CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D4PHI1Z2_CM_L5L6_L1D4PHI1Z2;
wire ME_L5L6_L1D4PHI1Z2_CM_L5L6_L1D4PHI1Z2_wr_en;
wire [5:0] CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI1Z2(
.data_in(ME_L5L6_L1D4PHI1Z2_CM_L5L6_L1D4PHI1Z2),
.enable(ME_L5L6_L1D4PHI1Z2_CM_L5L6_L1D4PHI1Z2_wr_en),
.number_out(CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D4PHI2Z1_CM_L5L6_L1D4PHI2Z1;
wire ME_L5L6_L1D4PHI2Z1_CM_L5L6_L1D4PHI2Z1_wr_en;
wire [5:0] CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI2Z1(
.data_in(ME_L5L6_L1D4PHI2Z1_CM_L5L6_L1D4PHI2Z1),
.enable(ME_L5L6_L1D4PHI2Z1_CM_L5L6_L1D4PHI2Z1_wr_en),
.number_out(CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D4PHI2Z2_CM_L5L6_L1D4PHI2Z2;
wire ME_L5L6_L1D4PHI2Z2_CM_L5L6_L1D4PHI2Z2_wr_en;
wire [5:0] CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI2Z2(
.data_in(ME_L5L6_L1D4PHI2Z2_CM_L5L6_L1D4PHI2Z2),
.enable(ME_L5L6_L1D4PHI2Z2_CM_L5L6_L1D4PHI2Z2_wr_en),
.number_out(CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D4PHI3Z1_CM_L5L6_L1D4PHI3Z1;
wire ME_L5L6_L1D4PHI3Z1_CM_L5L6_L1D4PHI3Z1_wr_en;
wire [5:0] CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI3Z1(
.data_in(ME_L5L6_L1D4PHI3Z1_CM_L5L6_L1D4PHI3Z1),
.enable(ME_L5L6_L1D4PHI3Z1_CM_L5L6_L1D4PHI3Z1_wr_en),
.number_out(CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L1D4PHI3Z2_CM_L5L6_L1D4PHI3Z2;
wire ME_L5L6_L1D4PHI3Z2_CM_L5L6_L1D4PHI3Z2_wr_en;
wire [5:0] CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI3Z2(
.data_in(ME_L5L6_L1D4PHI3Z2_CM_L5L6_L1D4PHI3Z2),
.enable(ME_L5L6_L1D4PHI3Z2_CM_L5L6_L1D4PHI3Z2_wr_en),
.number_out(CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L1D4_L5L6_AP_L5L6_L1D4;
wire PR_L1D4_L5L6_AP_L5L6_L1D4_wr_en;
wire [8:0] AP_L5L6_L1D4_MC_L5L6_L1D4_read_add;
wire [55:0] AP_L5L6_L1D4_MC_L5L6_L1D4;
AllProj #(1'b1) AP_L5L6_L1D4(
.data_in(PR_L1D4_L5L6_AP_L5L6_L1D4),
.enable(PR_L1D4_L5L6_AP_L5L6_L1D4_wr_en),
.read_add(AP_L5L6_L1D4_MC_L5L6_L1D4_read_add),
.data_out(AP_L5L6_L1D4_MC_L5L6_L1D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L1D4_AS_L1D4n3;
wire VMR_L1D4_AS_L1D4n3_wr_en;
wire [10:0] AS_L1D4n3_MC_L5L6_L1D4_read_add;
wire [35:0] AS_L1D4n3_MC_L5L6_L1D4;
AllStubs  AS_L1D4n3(
.data_in(VMR_L1D4_AS_L1D4n3),
.enable(VMR_L1D4_AS_L1D4n3_wr_en),
.read_add_MC(AS_L1D4n3_MC_L5L6_L1D4_read_add),
.data_out_MC(AS_L1D4n3_MC_L5L6_L1D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D3PHI1Z1_CM_L5L6_L2D3PHI1Z1;
wire ME_L5L6_L2D3PHI1Z1_CM_L5L6_L2D3PHI1Z1_wr_en;
wire [5:0] CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI1Z1(
.data_in(ME_L5L6_L2D3PHI1Z1_CM_L5L6_L2D3PHI1Z1),
.enable(ME_L5L6_L2D3PHI1Z1_CM_L5L6_L2D3PHI1Z1_wr_en),
.number_out(CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D3PHI1Z2_CM_L5L6_L2D3PHI1Z2;
wire ME_L5L6_L2D3PHI1Z2_CM_L5L6_L2D3PHI1Z2_wr_en;
wire [5:0] CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI1Z2(
.data_in(ME_L5L6_L2D3PHI1Z2_CM_L5L6_L2D3PHI1Z2),
.enable(ME_L5L6_L2D3PHI1Z2_CM_L5L6_L2D3PHI1Z2_wr_en),
.number_out(CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D3PHI2Z1_CM_L5L6_L2D3PHI2Z1;
wire ME_L5L6_L2D3PHI2Z1_CM_L5L6_L2D3PHI2Z1_wr_en;
wire [5:0] CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI2Z1(
.data_in(ME_L5L6_L2D3PHI2Z1_CM_L5L6_L2D3PHI2Z1),
.enable(ME_L5L6_L2D3PHI2Z1_CM_L5L6_L2D3PHI2Z1_wr_en),
.number_out(CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D3PHI2Z2_CM_L5L6_L2D3PHI2Z2;
wire ME_L5L6_L2D3PHI2Z2_CM_L5L6_L2D3PHI2Z2_wr_en;
wire [5:0] CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI2Z2(
.data_in(ME_L5L6_L2D3PHI2Z2_CM_L5L6_L2D3PHI2Z2),
.enable(ME_L5L6_L2D3PHI2Z2_CM_L5L6_L2D3PHI2Z2_wr_en),
.number_out(CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D3PHI3Z1_CM_L5L6_L2D3PHI3Z1;
wire ME_L5L6_L2D3PHI3Z1_CM_L5L6_L2D3PHI3Z1_wr_en;
wire [5:0] CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI3Z1(
.data_in(ME_L5L6_L2D3PHI3Z1_CM_L5L6_L2D3PHI3Z1),
.enable(ME_L5L6_L2D3PHI3Z1_CM_L5L6_L2D3PHI3Z1_wr_en),
.number_out(CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D3PHI3Z2_CM_L5L6_L2D3PHI3Z2;
wire ME_L5L6_L2D3PHI3Z2_CM_L5L6_L2D3PHI3Z2_wr_en;
wire [5:0] CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI3Z2(
.data_in(ME_L5L6_L2D3PHI3Z2_CM_L5L6_L2D3PHI3Z2),
.enable(ME_L5L6_L2D3PHI3Z2_CM_L5L6_L2D3PHI3Z2_wr_en),
.number_out(CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D3PHI4Z1_CM_L5L6_L2D3PHI4Z1;
wire ME_L5L6_L2D3PHI4Z1_CM_L5L6_L2D3PHI4Z1_wr_en;
wire [5:0] CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI4Z1(
.data_in(ME_L5L6_L2D3PHI4Z1_CM_L5L6_L2D3PHI4Z1),
.enable(ME_L5L6_L2D3PHI4Z1_CM_L5L6_L2D3PHI4Z1_wr_en),
.number_out(CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D3PHI4Z2_CM_L5L6_L2D3PHI4Z2;
wire ME_L5L6_L2D3PHI4Z2_CM_L5L6_L2D3PHI4Z2_wr_en;
wire [5:0] CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI4Z2(
.data_in(ME_L5L6_L2D3PHI4Z2_CM_L5L6_L2D3PHI4Z2),
.enable(ME_L5L6_L2D3PHI4Z2_CM_L5L6_L2D3PHI4Z2_wr_en),
.number_out(CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L2D3_L5L6_AP_L5L6_L2D3;
wire PR_L2D3_L5L6_AP_L5L6_L2D3_wr_en;
wire [8:0] AP_L5L6_L2D3_MC_L5L6_L2D3_read_add;
wire [55:0] AP_L5L6_L2D3_MC_L5L6_L2D3;
AllProj #(1'b1) AP_L5L6_L2D3(
.data_in(PR_L2D3_L5L6_AP_L5L6_L2D3),
.enable(PR_L2D3_L5L6_AP_L5L6_L2D3_wr_en),
.read_add(AP_L5L6_L2D3_MC_L5L6_L2D3_read_add),
.data_out(AP_L5L6_L2D3_MC_L5L6_L2D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L2D3_AS_L2D3n3;
wire VMR_L2D3_AS_L2D3n3_wr_en;
wire [10:0] AS_L2D3n3_MC_L5L6_L2D3_read_add;
wire [35:0] AS_L2D3n3_MC_L5L6_L2D3;
AllStubs  AS_L2D3n3(
.data_in(VMR_L2D3_AS_L2D3n3),
.enable(VMR_L2D3_AS_L2D3n3_wr_en),
.read_add_MC(AS_L2D3n3_MC_L5L6_L2D3_read_add),
.data_out_MC(AS_L2D3n3_MC_L5L6_L2D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D4PHI1Z1_CM_L5L6_L2D4PHI1Z1;
wire ME_L5L6_L2D4PHI1Z1_CM_L5L6_L2D4PHI1Z1_wr_en;
wire [5:0] CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI1Z1(
.data_in(ME_L5L6_L2D4PHI1Z1_CM_L5L6_L2D4PHI1Z1),
.enable(ME_L5L6_L2D4PHI1Z1_CM_L5L6_L2D4PHI1Z1_wr_en),
.number_out(CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D4PHI1Z2_CM_L5L6_L2D4PHI1Z2;
wire ME_L5L6_L2D4PHI1Z2_CM_L5L6_L2D4PHI1Z2_wr_en;
wire [5:0] CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI1Z2(
.data_in(ME_L5L6_L2D4PHI1Z2_CM_L5L6_L2D4PHI1Z2),
.enable(ME_L5L6_L2D4PHI1Z2_CM_L5L6_L2D4PHI1Z2_wr_en),
.number_out(CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D4PHI2Z1_CM_L5L6_L2D4PHI2Z1;
wire ME_L5L6_L2D4PHI2Z1_CM_L5L6_L2D4PHI2Z1_wr_en;
wire [5:0] CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI2Z1(
.data_in(ME_L5L6_L2D4PHI2Z1_CM_L5L6_L2D4PHI2Z1),
.enable(ME_L5L6_L2D4PHI2Z1_CM_L5L6_L2D4PHI2Z1_wr_en),
.number_out(CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D4PHI2Z2_CM_L5L6_L2D4PHI2Z2;
wire ME_L5L6_L2D4PHI2Z2_CM_L5L6_L2D4PHI2Z2_wr_en;
wire [5:0] CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI2Z2(
.data_in(ME_L5L6_L2D4PHI2Z2_CM_L5L6_L2D4PHI2Z2),
.enable(ME_L5L6_L2D4PHI2Z2_CM_L5L6_L2D4PHI2Z2_wr_en),
.number_out(CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D4PHI3Z1_CM_L5L6_L2D4PHI3Z1;
wire ME_L5L6_L2D4PHI3Z1_CM_L5L6_L2D4PHI3Z1_wr_en;
wire [5:0] CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI3Z1(
.data_in(ME_L5L6_L2D4PHI3Z1_CM_L5L6_L2D4PHI3Z1),
.enable(ME_L5L6_L2D4PHI3Z1_CM_L5L6_L2D4PHI3Z1_wr_en),
.number_out(CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D4PHI3Z2_CM_L5L6_L2D4PHI3Z2;
wire ME_L5L6_L2D4PHI3Z2_CM_L5L6_L2D4PHI3Z2_wr_en;
wire [5:0] CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI3Z2(
.data_in(ME_L5L6_L2D4PHI3Z2_CM_L5L6_L2D4PHI3Z2),
.enable(ME_L5L6_L2D4PHI3Z2_CM_L5L6_L2D4PHI3Z2_wr_en),
.number_out(CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D4PHI4Z1_CM_L5L6_L2D4PHI4Z1;
wire ME_L5L6_L2D4PHI4Z1_CM_L5L6_L2D4PHI4Z1_wr_en;
wire [5:0] CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI4Z1(
.data_in(ME_L5L6_L2D4PHI4Z1_CM_L5L6_L2D4PHI4Z1),
.enable(ME_L5L6_L2D4PHI4Z1_CM_L5L6_L2D4PHI4Z1_wr_en),
.number_out(CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L2D4PHI4Z2_CM_L5L6_L2D4PHI4Z2;
wire ME_L5L6_L2D4PHI4Z2_CM_L5L6_L2D4PHI4Z2_wr_en;
wire [5:0] CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI4Z2(
.data_in(ME_L5L6_L2D4PHI4Z2_CM_L5L6_L2D4PHI4Z2),
.enable(ME_L5L6_L2D4PHI4Z2_CM_L5L6_L2D4PHI4Z2_wr_en),
.number_out(CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L2D4_L5L6_AP_L5L6_L2D4;
wire PR_L2D4_L5L6_AP_L5L6_L2D4_wr_en;
wire [8:0] AP_L5L6_L2D4_MC_L5L6_L2D4_read_add;
wire [55:0] AP_L5L6_L2D4_MC_L5L6_L2D4;
AllProj #(1'b1) AP_L5L6_L2D4(
.data_in(PR_L2D4_L5L6_AP_L5L6_L2D4),
.enable(PR_L2D4_L5L6_AP_L5L6_L2D4_wr_en),
.read_add(AP_L5L6_L2D4_MC_L5L6_L2D4_read_add),
.data_out(AP_L5L6_L2D4_MC_L5L6_L2D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L2D4_AS_L2D4n4;
wire VMR_L2D4_AS_L2D4n4_wr_en;
wire [10:0] AS_L2D4n4_MC_L5L6_L2D4_read_add;
wire [35:0] AS_L2D4n4_MC_L5L6_L2D4;
AllStubs  AS_L2D4n4(
.data_in(VMR_L2D4_AS_L2D4n4),
.enable(VMR_L2D4_AS_L2D4n4_wr_en),
.read_add_MC(AS_L2D4n4_MC_L5L6_L2D4_read_add),
.data_out_MC(AS_L2D4n4_MC_L5L6_L2D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D3PHI1Z1_CM_L5L6_L3D3PHI1Z1;
wire ME_L5L6_L3D3PHI1Z1_CM_L5L6_L3D3PHI1Z1_wr_en;
wire [5:0] CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI1Z1(
.data_in(ME_L5L6_L3D3PHI1Z1_CM_L5L6_L3D3PHI1Z1),
.enable(ME_L5L6_L3D3PHI1Z1_CM_L5L6_L3D3PHI1Z1_wr_en),
.number_out(CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D3PHI1Z2_CM_L5L6_L3D3PHI1Z2;
wire ME_L5L6_L3D3PHI1Z2_CM_L5L6_L3D3PHI1Z2_wr_en;
wire [5:0] CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI1Z2(
.data_in(ME_L5L6_L3D3PHI1Z2_CM_L5L6_L3D3PHI1Z2),
.enable(ME_L5L6_L3D3PHI1Z2_CM_L5L6_L3D3PHI1Z2_wr_en),
.number_out(CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D3PHI2Z1_CM_L5L6_L3D3PHI2Z1;
wire ME_L5L6_L3D3PHI2Z1_CM_L5L6_L3D3PHI2Z1_wr_en;
wire [5:0] CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI2Z1(
.data_in(ME_L5L6_L3D3PHI2Z1_CM_L5L6_L3D3PHI2Z1),
.enable(ME_L5L6_L3D3PHI2Z1_CM_L5L6_L3D3PHI2Z1_wr_en),
.number_out(CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D3PHI2Z2_CM_L5L6_L3D3PHI2Z2;
wire ME_L5L6_L3D3PHI2Z2_CM_L5L6_L3D3PHI2Z2_wr_en;
wire [5:0] CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI2Z2(
.data_in(ME_L5L6_L3D3PHI2Z2_CM_L5L6_L3D3PHI2Z2),
.enable(ME_L5L6_L3D3PHI2Z2_CM_L5L6_L3D3PHI2Z2_wr_en),
.number_out(CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D3PHI3Z1_CM_L5L6_L3D3PHI3Z1;
wire ME_L5L6_L3D3PHI3Z1_CM_L5L6_L3D3PHI3Z1_wr_en;
wire [5:0] CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI3Z1(
.data_in(ME_L5L6_L3D3PHI3Z1_CM_L5L6_L3D3PHI3Z1),
.enable(ME_L5L6_L3D3PHI3Z1_CM_L5L6_L3D3PHI3Z1_wr_en),
.number_out(CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D3PHI3Z2_CM_L5L6_L3D3PHI3Z2;
wire ME_L5L6_L3D3PHI3Z2_CM_L5L6_L3D3PHI3Z2_wr_en;
wire [5:0] CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI3Z2(
.data_in(ME_L5L6_L3D3PHI3Z2_CM_L5L6_L3D3PHI3Z2),
.enable(ME_L5L6_L3D3PHI3Z2_CM_L5L6_L3D3PHI3Z2_wr_en),
.number_out(CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L3D3_L5L6_AP_L5L6_L3D3;
wire PR_L3D3_L5L6_AP_L5L6_L3D3_wr_en;
wire [8:0] AP_L5L6_L3D3_MC_L5L6_L3D3_read_add;
wire [55:0] AP_L5L6_L3D3_MC_L5L6_L3D3;
AllProj #(1'b1) AP_L5L6_L3D3(
.data_in(PR_L3D3_L5L6_AP_L5L6_L3D3),
.enable(PR_L3D3_L5L6_AP_L5L6_L3D3_wr_en),
.read_add(AP_L5L6_L3D3_MC_L5L6_L3D3_read_add),
.data_out(AP_L5L6_L3D3_MC_L5L6_L3D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L3D3_AS_L3D3n3;
wire VMR_L3D3_AS_L3D3n3_wr_en;
wire [10:0] AS_L3D3n3_MC_L5L6_L3D3_read_add;
wire [35:0] AS_L3D3n3_MC_L5L6_L3D3;
AllStubs  AS_L3D3n3(
.data_in(VMR_L3D3_AS_L3D3n3),
.enable(VMR_L3D3_AS_L3D3n3_wr_en),
.read_add_MC(AS_L3D3n3_MC_L5L6_L3D3_read_add),
.data_out_MC(AS_L3D3n3_MC_L5L6_L3D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D4PHI1Z1_CM_L5L6_L3D4PHI1Z1;
wire ME_L5L6_L3D4PHI1Z1_CM_L5L6_L3D4PHI1Z1_wr_en;
wire [5:0] CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI1Z1(
.data_in(ME_L5L6_L3D4PHI1Z1_CM_L5L6_L3D4PHI1Z1),
.enable(ME_L5L6_L3D4PHI1Z1_CM_L5L6_L3D4PHI1Z1_wr_en),
.number_out(CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D4PHI1Z2_CM_L5L6_L3D4PHI1Z2;
wire ME_L5L6_L3D4PHI1Z2_CM_L5L6_L3D4PHI1Z2_wr_en;
wire [5:0] CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI1Z2(
.data_in(ME_L5L6_L3D4PHI1Z2_CM_L5L6_L3D4PHI1Z2),
.enable(ME_L5L6_L3D4PHI1Z2_CM_L5L6_L3D4PHI1Z2_wr_en),
.number_out(CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D4PHI2Z1_CM_L5L6_L3D4PHI2Z1;
wire ME_L5L6_L3D4PHI2Z1_CM_L5L6_L3D4PHI2Z1_wr_en;
wire [5:0] CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI2Z1(
.data_in(ME_L5L6_L3D4PHI2Z1_CM_L5L6_L3D4PHI2Z1),
.enable(ME_L5L6_L3D4PHI2Z1_CM_L5L6_L3D4PHI2Z1_wr_en),
.number_out(CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D4PHI2Z2_CM_L5L6_L3D4PHI2Z2;
wire ME_L5L6_L3D4PHI2Z2_CM_L5L6_L3D4PHI2Z2_wr_en;
wire [5:0] CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI2Z2(
.data_in(ME_L5L6_L3D4PHI2Z2_CM_L5L6_L3D4PHI2Z2),
.enable(ME_L5L6_L3D4PHI2Z2_CM_L5L6_L3D4PHI2Z2_wr_en),
.number_out(CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D4PHI3Z1_CM_L5L6_L3D4PHI3Z1;
wire ME_L5L6_L3D4PHI3Z1_CM_L5L6_L3D4PHI3Z1_wr_en;
wire [5:0] CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI3Z1(
.data_in(ME_L5L6_L3D4PHI3Z1_CM_L5L6_L3D4PHI3Z1),
.enable(ME_L5L6_L3D4PHI3Z1_CM_L5L6_L3D4PHI3Z1_wr_en),
.number_out(CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L3D4PHI3Z2_CM_L5L6_L3D4PHI3Z2;
wire ME_L5L6_L3D4PHI3Z2_CM_L5L6_L3D4PHI3Z2_wr_en;
wire [5:0] CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI3Z2(
.data_in(ME_L5L6_L3D4PHI3Z2_CM_L5L6_L3D4PHI3Z2),
.enable(ME_L5L6_L3D4PHI3Z2_CM_L5L6_L3D4PHI3Z2_wr_en),
.number_out(CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L3D4_L5L6_AP_L5L6_L3D4;
wire PR_L3D4_L5L6_AP_L5L6_L3D4_wr_en;
wire [8:0] AP_L5L6_L3D4_MC_L5L6_L3D4_read_add;
wire [55:0] AP_L5L6_L3D4_MC_L5L6_L3D4;
AllProj #(1'b1) AP_L5L6_L3D4(
.data_in(PR_L3D4_L5L6_AP_L5L6_L3D4),
.enable(PR_L3D4_L5L6_AP_L5L6_L3D4_wr_en),
.read_add(AP_L5L6_L3D4_MC_L5L6_L3D4_read_add),
.data_out(AP_L5L6_L3D4_MC_L5L6_L3D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L3D4_AS_L3D4n2;
wire VMR_L3D4_AS_L3D4n2_wr_en;
wire [10:0] AS_L3D4n2_MC_L5L6_L3D4_read_add;
wire [35:0] AS_L3D4n2_MC_L5L6_L3D4;
AllStubs  AS_L3D4n2(
.data_in(VMR_L3D4_AS_L3D4n2),
.enable(VMR_L3D4_AS_L3D4n2_wr_en),
.read_add_MC(AS_L3D4n2_MC_L5L6_L3D4_read_add),
.data_out_MC(AS_L3D4n2_MC_L5L6_L3D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D3PHI1Z1_CM_L5L6_L4D3PHI1Z1;
wire ME_L5L6_L4D3PHI1Z1_CM_L5L6_L4D3PHI1Z1_wr_en;
wire [5:0] CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI1Z1(
.data_in(ME_L5L6_L4D3PHI1Z1_CM_L5L6_L4D3PHI1Z1),
.enable(ME_L5L6_L4D3PHI1Z1_CM_L5L6_L4D3PHI1Z1_wr_en),
.number_out(CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D3PHI1Z2_CM_L5L6_L4D3PHI1Z2;
wire ME_L5L6_L4D3PHI1Z2_CM_L5L6_L4D3PHI1Z2_wr_en;
wire [5:0] CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI1Z2(
.data_in(ME_L5L6_L4D3PHI1Z2_CM_L5L6_L4D3PHI1Z2),
.enable(ME_L5L6_L4D3PHI1Z2_CM_L5L6_L4D3PHI1Z2_wr_en),
.number_out(CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D3PHI2Z1_CM_L5L6_L4D3PHI2Z1;
wire ME_L5L6_L4D3PHI2Z1_CM_L5L6_L4D3PHI2Z1_wr_en;
wire [5:0] CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI2Z1(
.data_in(ME_L5L6_L4D3PHI2Z1_CM_L5L6_L4D3PHI2Z1),
.enable(ME_L5L6_L4D3PHI2Z1_CM_L5L6_L4D3PHI2Z1_wr_en),
.number_out(CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D3PHI2Z2_CM_L5L6_L4D3PHI2Z2;
wire ME_L5L6_L4D3PHI2Z2_CM_L5L6_L4D3PHI2Z2_wr_en;
wire [5:0] CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI2Z2(
.data_in(ME_L5L6_L4D3PHI2Z2_CM_L5L6_L4D3PHI2Z2),
.enable(ME_L5L6_L4D3PHI2Z2_CM_L5L6_L4D3PHI2Z2_wr_en),
.number_out(CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D3PHI3Z1_CM_L5L6_L4D3PHI3Z1;
wire ME_L5L6_L4D3PHI3Z1_CM_L5L6_L4D3PHI3Z1_wr_en;
wire [5:0] CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI3Z1(
.data_in(ME_L5L6_L4D3PHI3Z1_CM_L5L6_L4D3PHI3Z1),
.enable(ME_L5L6_L4D3PHI3Z1_CM_L5L6_L4D3PHI3Z1_wr_en),
.number_out(CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D3PHI3Z2_CM_L5L6_L4D3PHI3Z2;
wire ME_L5L6_L4D3PHI3Z2_CM_L5L6_L4D3PHI3Z2_wr_en;
wire [5:0] CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI3Z2(
.data_in(ME_L5L6_L4D3PHI3Z2_CM_L5L6_L4D3PHI3Z2),
.enable(ME_L5L6_L4D3PHI3Z2_CM_L5L6_L4D3PHI3Z2_wr_en),
.number_out(CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D3PHI4Z1_CM_L5L6_L4D3PHI4Z1;
wire ME_L5L6_L4D3PHI4Z1_CM_L5L6_L4D3PHI4Z1_wr_en;
wire [5:0] CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI4Z1(
.data_in(ME_L5L6_L4D3PHI4Z1_CM_L5L6_L4D3PHI4Z1),
.enable(ME_L5L6_L4D3PHI4Z1_CM_L5L6_L4D3PHI4Z1_wr_en),
.number_out(CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D3PHI4Z2_CM_L5L6_L4D3PHI4Z2;
wire ME_L5L6_L4D3PHI4Z2_CM_L5L6_L4D3PHI4Z2_wr_en;
wire [5:0] CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI4Z2(
.data_in(ME_L5L6_L4D3PHI4Z2_CM_L5L6_L4D3PHI4Z2),
.enable(ME_L5L6_L4D3PHI4Z2_CM_L5L6_L4D3PHI4Z2_wr_en),
.number_out(CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L4D3_L5L6_AP_L5L6_L4D3;
wire PR_L4D3_L5L6_AP_L5L6_L4D3_wr_en;
wire [8:0] AP_L5L6_L4D3_MC_L5L6_L4D3_read_add;
wire [55:0] AP_L5L6_L4D3_MC_L5L6_L4D3;
AllProj #(1'b0) AP_L5L6_L4D3(
.data_in(PR_L4D3_L5L6_AP_L5L6_L4D3),
.enable(PR_L4D3_L5L6_AP_L5L6_L4D3_wr_en),
.read_add(AP_L5L6_L4D3_MC_L5L6_L4D3_read_add),
.data_out(AP_L5L6_L4D3_MC_L5L6_L4D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L4D3_AS_L4D3n2;
wire VMR_L4D3_AS_L4D3n2_wr_en;
wire [10:0] AS_L4D3n2_MC_L5L6_L4D3_read_add;
wire [35:0] AS_L4D3n2_MC_L5L6_L4D3;
AllStubs  AS_L4D3n2(
.data_in(VMR_L4D3_AS_L4D3n2),
.enable(VMR_L4D3_AS_L4D3n2_wr_en),
.read_add_MC(AS_L4D3n2_MC_L5L6_L4D3_read_add),
.data_out_MC(AS_L4D3n2_MC_L5L6_L4D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D4PHI1Z1_CM_L5L6_L4D4PHI1Z1;
wire ME_L5L6_L4D4PHI1Z1_CM_L5L6_L4D4PHI1Z1_wr_en;
wire [5:0] CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI1Z1(
.data_in(ME_L5L6_L4D4PHI1Z1_CM_L5L6_L4D4PHI1Z1),
.enable(ME_L5L6_L4D4PHI1Z1_CM_L5L6_L4D4PHI1Z1_wr_en),
.number_out(CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D4PHI1Z2_CM_L5L6_L4D4PHI1Z2;
wire ME_L5L6_L4D4PHI1Z2_CM_L5L6_L4D4PHI1Z2_wr_en;
wire [5:0] CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI1Z2(
.data_in(ME_L5L6_L4D4PHI1Z2_CM_L5L6_L4D4PHI1Z2),
.enable(ME_L5L6_L4D4PHI1Z2_CM_L5L6_L4D4PHI1Z2_wr_en),
.number_out(CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D4PHI2Z1_CM_L5L6_L4D4PHI2Z1;
wire ME_L5L6_L4D4PHI2Z1_CM_L5L6_L4D4PHI2Z1_wr_en;
wire [5:0] CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI2Z1(
.data_in(ME_L5L6_L4D4PHI2Z1_CM_L5L6_L4D4PHI2Z1),
.enable(ME_L5L6_L4D4PHI2Z1_CM_L5L6_L4D4PHI2Z1_wr_en),
.number_out(CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D4PHI2Z2_CM_L5L6_L4D4PHI2Z2;
wire ME_L5L6_L4D4PHI2Z2_CM_L5L6_L4D4PHI2Z2_wr_en;
wire [5:0] CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI2Z2(
.data_in(ME_L5L6_L4D4PHI2Z2_CM_L5L6_L4D4PHI2Z2),
.enable(ME_L5L6_L4D4PHI2Z2_CM_L5L6_L4D4PHI2Z2_wr_en),
.number_out(CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D4PHI3Z1_CM_L5L6_L4D4PHI3Z1;
wire ME_L5L6_L4D4PHI3Z1_CM_L5L6_L4D4PHI3Z1_wr_en;
wire [5:0] CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI3Z1(
.data_in(ME_L5L6_L4D4PHI3Z1_CM_L5L6_L4D4PHI3Z1),
.enable(ME_L5L6_L4D4PHI3Z1_CM_L5L6_L4D4PHI3Z1_wr_en),
.number_out(CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D4PHI3Z2_CM_L5L6_L4D4PHI3Z2;
wire ME_L5L6_L4D4PHI3Z2_CM_L5L6_L4D4PHI3Z2_wr_en;
wire [5:0] CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI3Z2(
.data_in(ME_L5L6_L4D4PHI3Z2_CM_L5L6_L4D4PHI3Z2),
.enable(ME_L5L6_L4D4PHI3Z2_CM_L5L6_L4D4PHI3Z2_wr_en),
.number_out(CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D4PHI4Z1_CM_L5L6_L4D4PHI4Z1;
wire ME_L5L6_L4D4PHI4Z1_CM_L5L6_L4D4PHI4Z1_wr_en;
wire [5:0] CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI4Z1(
.data_in(ME_L5L6_L4D4PHI4Z1_CM_L5L6_L4D4PHI4Z1),
.enable(ME_L5L6_L4D4PHI4Z1_CM_L5L6_L4D4PHI4Z1_wr_en),
.number_out(CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L5L6_L4D4PHI4Z2_CM_L5L6_L4D4PHI4Z2;
wire ME_L5L6_L4D4PHI4Z2_CM_L5L6_L4D4PHI4Z2_wr_en;
wire [5:0] CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI4Z2(
.data_in(ME_L5L6_L4D4PHI4Z2_CM_L5L6_L4D4PHI4Z2),
.enable(ME_L5L6_L4D4PHI4Z2_CM_L5L6_L4D4PHI4Z2_wr_en),
.number_out(CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L4D4_L5L6_AP_L5L6_L4D4;
wire PR_L4D4_L5L6_AP_L5L6_L4D4_wr_en;
wire [8:0] AP_L5L6_L4D4_MC_L5L6_L4D4_read_add;
wire [55:0] AP_L5L6_L4D4_MC_L5L6_L4D4;
AllProj #(1'b0) AP_L5L6_L4D4(
.data_in(PR_L4D4_L5L6_AP_L5L6_L4D4),
.enable(PR_L4D4_L5L6_AP_L5L6_L4D4_wr_en),
.read_add(AP_L5L6_L4D4_MC_L5L6_L4D4_read_add),
.data_out(AP_L5L6_L4D4_MC_L5L6_L4D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L4D4_AS_L4D4n3;
wire VMR_L4D4_AS_L4D4n3_wr_en;
wire [10:0] AS_L4D4n3_MC_L5L6_L4D4_read_add;
wire [35:0] AS_L4D4n3_MC_L5L6_L4D4;
AllStubs  AS_L4D4n3(
.data_in(VMR_L4D4_AS_L4D4n3),
.enable(VMR_L4D4_AS_L4D4n3_wr_en),
.read_add_MC(AS_L4D4n3_MC_L5L6_L4D4_read_add),
.data_out_MC(AS_L4D4n3_MC_L5L6_L4D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D3PHI1Z1_CM_L1L2_L3D3PHI1Z1;
wire ME_L1L2_L3D3PHI1Z1_CM_L1L2_L3D3PHI1Z1_wr_en;
wire [5:0] CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI1Z1(
.data_in(ME_L1L2_L3D3PHI1Z1_CM_L1L2_L3D3PHI1Z1),
.enable(ME_L1L2_L3D3PHI1Z1_CM_L1L2_L3D3PHI1Z1_wr_en),
.number_out(CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D3PHI1Z2_CM_L1L2_L3D3PHI1Z2;
wire ME_L1L2_L3D3PHI1Z2_CM_L1L2_L3D3PHI1Z2_wr_en;
wire [5:0] CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI1Z2(
.data_in(ME_L1L2_L3D3PHI1Z2_CM_L1L2_L3D3PHI1Z2),
.enable(ME_L1L2_L3D3PHI1Z2_CM_L1L2_L3D3PHI1Z2_wr_en),
.number_out(CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D3PHI2Z1_CM_L1L2_L3D3PHI2Z1;
wire ME_L1L2_L3D3PHI2Z1_CM_L1L2_L3D3PHI2Z1_wr_en;
wire [5:0] CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI2Z1(
.data_in(ME_L1L2_L3D3PHI2Z1_CM_L1L2_L3D3PHI2Z1),
.enable(ME_L1L2_L3D3PHI2Z1_CM_L1L2_L3D3PHI2Z1_wr_en),
.number_out(CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D3PHI2Z2_CM_L1L2_L3D3PHI2Z2;
wire ME_L1L2_L3D3PHI2Z2_CM_L1L2_L3D3PHI2Z2_wr_en;
wire [5:0] CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI2Z2(
.data_in(ME_L1L2_L3D3PHI2Z2_CM_L1L2_L3D3PHI2Z2),
.enable(ME_L1L2_L3D3PHI2Z2_CM_L1L2_L3D3PHI2Z2_wr_en),
.number_out(CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D3PHI3Z1_CM_L1L2_L3D3PHI3Z1;
wire ME_L1L2_L3D3PHI3Z1_CM_L1L2_L3D3PHI3Z1_wr_en;
wire [5:0] CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI3Z1(
.data_in(ME_L1L2_L3D3PHI3Z1_CM_L1L2_L3D3PHI3Z1),
.enable(ME_L1L2_L3D3PHI3Z1_CM_L1L2_L3D3PHI3Z1_wr_en),
.number_out(CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D3PHI3Z2_CM_L1L2_L3D3PHI3Z2;
wire ME_L1L2_L3D3PHI3Z2_CM_L1L2_L3D3PHI3Z2_wr_en;
wire [5:0] CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI3Z2(
.data_in(ME_L1L2_L3D3PHI3Z2_CM_L1L2_L3D3PHI3Z2),
.enable(ME_L1L2_L3D3PHI3Z2_CM_L1L2_L3D3PHI3Z2_wr_en),
.number_out(CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L3D3_L1L2_AP_L1L2_L3D3;
wire PR_L3D3_L1L2_AP_L1L2_L3D3_wr_en;
wire [8:0] AP_L1L2_L3D3_MC_L1L2_L3D3_read_add;
wire [55:0] AP_L1L2_L3D3_MC_L1L2_L3D3;
AllProj #(1'b1) AP_L1L2_L3D3(
.data_in(PR_L3D3_L1L2_AP_L1L2_L3D3),
.enable(PR_L3D3_L1L2_AP_L1L2_L3D3_wr_en),
.read_add(AP_L1L2_L3D3_MC_L1L2_L3D3_read_add),
.data_out(AP_L1L2_L3D3_MC_L1L2_L3D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L3D3_AS_L3D3n4;
wire VMR_L3D3_AS_L3D3n4_wr_en;
wire [10:0] AS_L3D3n4_MC_L1L2_L3D3_read_add;
wire [35:0] AS_L3D3n4_MC_L1L2_L3D3;
AllStubs  AS_L3D3n4(
.data_in(VMR_L3D3_AS_L3D3n4),
.enable(VMR_L3D3_AS_L3D3n4_wr_en),
.read_add_MC(AS_L3D3n4_MC_L1L2_L3D3_read_add),
.data_out_MC(AS_L3D3n4_MC_L1L2_L3D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D4PHI1Z1_CM_L1L2_L3D4PHI1Z1;
wire ME_L1L2_L3D4PHI1Z1_CM_L1L2_L3D4PHI1Z1_wr_en;
wire [5:0] CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI1Z1(
.data_in(ME_L1L2_L3D4PHI1Z1_CM_L1L2_L3D4PHI1Z1),
.enable(ME_L1L2_L3D4PHI1Z1_CM_L1L2_L3D4PHI1Z1_wr_en),
.number_out(CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D4PHI1Z2_CM_L1L2_L3D4PHI1Z2;
wire ME_L1L2_L3D4PHI1Z2_CM_L1L2_L3D4PHI1Z2_wr_en;
wire [5:0] CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI1Z2(
.data_in(ME_L1L2_L3D4PHI1Z2_CM_L1L2_L3D4PHI1Z2),
.enable(ME_L1L2_L3D4PHI1Z2_CM_L1L2_L3D4PHI1Z2_wr_en),
.number_out(CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D4PHI2Z1_CM_L1L2_L3D4PHI2Z1;
wire ME_L1L2_L3D4PHI2Z1_CM_L1L2_L3D4PHI2Z1_wr_en;
wire [5:0] CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI2Z1(
.data_in(ME_L1L2_L3D4PHI2Z1_CM_L1L2_L3D4PHI2Z1),
.enable(ME_L1L2_L3D4PHI2Z1_CM_L1L2_L3D4PHI2Z1_wr_en),
.number_out(CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D4PHI2Z2_CM_L1L2_L3D4PHI2Z2;
wire ME_L1L2_L3D4PHI2Z2_CM_L1L2_L3D4PHI2Z2_wr_en;
wire [5:0] CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI2Z2(
.data_in(ME_L1L2_L3D4PHI2Z2_CM_L1L2_L3D4PHI2Z2),
.enable(ME_L1L2_L3D4PHI2Z2_CM_L1L2_L3D4PHI2Z2_wr_en),
.number_out(CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D4PHI3Z1_CM_L1L2_L3D4PHI3Z1;
wire ME_L1L2_L3D4PHI3Z1_CM_L1L2_L3D4PHI3Z1_wr_en;
wire [5:0] CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI3Z1(
.data_in(ME_L1L2_L3D4PHI3Z1_CM_L1L2_L3D4PHI3Z1),
.enable(ME_L1L2_L3D4PHI3Z1_CM_L1L2_L3D4PHI3Z1_wr_en),
.number_out(CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L3D4PHI3Z2_CM_L1L2_L3D4PHI3Z2;
wire ME_L1L2_L3D4PHI3Z2_CM_L1L2_L3D4PHI3Z2_wr_en;
wire [5:0] CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI3Z2(
.data_in(ME_L1L2_L3D4PHI3Z2_CM_L1L2_L3D4PHI3Z2),
.enable(ME_L1L2_L3D4PHI3Z2_CM_L1L2_L3D4PHI3Z2_wr_en),
.number_out(CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L3D4_L1L2_AP_L1L2_L3D4;
wire PR_L3D4_L1L2_AP_L1L2_L3D4_wr_en;
wire [8:0] AP_L1L2_L3D4_MC_L1L2_L3D4_read_add;
wire [55:0] AP_L1L2_L3D4_MC_L1L2_L3D4;
AllProj #(1'b1) AP_L1L2_L3D4(
.data_in(PR_L3D4_L1L2_AP_L1L2_L3D4),
.enable(PR_L3D4_L1L2_AP_L1L2_L3D4_wr_en),
.read_add(AP_L1L2_L3D4_MC_L1L2_L3D4_read_add),
.data_out(AP_L1L2_L3D4_MC_L1L2_L3D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L3D4_AS_L3D4n3;
wire VMR_L3D4_AS_L3D4n3_wr_en;
wire [10:0] AS_L3D4n3_MC_L1L2_L3D4_read_add;
wire [35:0] AS_L3D4n3_MC_L1L2_L3D4;
AllStubs  AS_L3D4n3(
.data_in(VMR_L3D4_AS_L3D4n3),
.enable(VMR_L3D4_AS_L3D4n3_wr_en),
.read_add_MC(AS_L3D4n3_MC_L1L2_L3D4_read_add),
.data_out_MC(AS_L3D4n3_MC_L1L2_L3D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D3PHI1Z1_CM_L1L2_L4D3PHI1Z1;
wire ME_L1L2_L4D3PHI1Z1_CM_L1L2_L4D3PHI1Z1_wr_en;
wire [5:0] CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI1Z1(
.data_in(ME_L1L2_L4D3PHI1Z1_CM_L1L2_L4D3PHI1Z1),
.enable(ME_L1L2_L4D3PHI1Z1_CM_L1L2_L4D3PHI1Z1_wr_en),
.number_out(CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D3PHI1Z2_CM_L1L2_L4D3PHI1Z2;
wire ME_L1L2_L4D3PHI1Z2_CM_L1L2_L4D3PHI1Z2_wr_en;
wire [5:0] CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI1Z2(
.data_in(ME_L1L2_L4D3PHI1Z2_CM_L1L2_L4D3PHI1Z2),
.enable(ME_L1L2_L4D3PHI1Z2_CM_L1L2_L4D3PHI1Z2_wr_en),
.number_out(CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D3PHI2Z1_CM_L1L2_L4D3PHI2Z1;
wire ME_L1L2_L4D3PHI2Z1_CM_L1L2_L4D3PHI2Z1_wr_en;
wire [5:0] CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI2Z1(
.data_in(ME_L1L2_L4D3PHI2Z1_CM_L1L2_L4D3PHI2Z1),
.enable(ME_L1L2_L4D3PHI2Z1_CM_L1L2_L4D3PHI2Z1_wr_en),
.number_out(CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D3PHI2Z2_CM_L1L2_L4D3PHI2Z2;
wire ME_L1L2_L4D3PHI2Z2_CM_L1L2_L4D3PHI2Z2_wr_en;
wire [5:0] CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI2Z2(
.data_in(ME_L1L2_L4D3PHI2Z2_CM_L1L2_L4D3PHI2Z2),
.enable(ME_L1L2_L4D3PHI2Z2_CM_L1L2_L4D3PHI2Z2_wr_en),
.number_out(CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D3PHI3Z1_CM_L1L2_L4D3PHI3Z1;
wire ME_L1L2_L4D3PHI3Z1_CM_L1L2_L4D3PHI3Z1_wr_en;
wire [5:0] CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI3Z1(
.data_in(ME_L1L2_L4D3PHI3Z1_CM_L1L2_L4D3PHI3Z1),
.enable(ME_L1L2_L4D3PHI3Z1_CM_L1L2_L4D3PHI3Z1_wr_en),
.number_out(CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D3PHI3Z2_CM_L1L2_L4D3PHI3Z2;
wire ME_L1L2_L4D3PHI3Z2_CM_L1L2_L4D3PHI3Z2_wr_en;
wire [5:0] CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI3Z2(
.data_in(ME_L1L2_L4D3PHI3Z2_CM_L1L2_L4D3PHI3Z2),
.enable(ME_L1L2_L4D3PHI3Z2_CM_L1L2_L4D3PHI3Z2_wr_en),
.number_out(CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D3PHI4Z1_CM_L1L2_L4D3PHI4Z1;
wire ME_L1L2_L4D3PHI4Z1_CM_L1L2_L4D3PHI4Z1_wr_en;
wire [5:0] CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI4Z1(
.data_in(ME_L1L2_L4D3PHI4Z1_CM_L1L2_L4D3PHI4Z1),
.enable(ME_L1L2_L4D3PHI4Z1_CM_L1L2_L4D3PHI4Z1_wr_en),
.number_out(CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D3PHI4Z2_CM_L1L2_L4D3PHI4Z2;
wire ME_L1L2_L4D3PHI4Z2_CM_L1L2_L4D3PHI4Z2_wr_en;
wire [5:0] CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI4Z2(
.data_in(ME_L1L2_L4D3PHI4Z2_CM_L1L2_L4D3PHI4Z2),
.enable(ME_L1L2_L4D3PHI4Z2_CM_L1L2_L4D3PHI4Z2_wr_en),
.number_out(CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L4D3_L1L2_AP_L1L2_L4D3;
wire PR_L4D3_L1L2_AP_L1L2_L4D3_wr_en;
wire [8:0] AP_L1L2_L4D3_MC_L1L2_L4D3_read_add;
wire [55:0] AP_L1L2_L4D3_MC_L1L2_L4D3;
AllProj #(1'b0) AP_L1L2_L4D3(
.data_in(PR_L4D3_L1L2_AP_L1L2_L4D3),
.enable(PR_L4D3_L1L2_AP_L1L2_L4D3_wr_en),
.read_add(AP_L1L2_L4D3_MC_L1L2_L4D3_read_add),
.data_out(AP_L1L2_L4D3_MC_L1L2_L4D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L4D3_AS_L4D3n3;
wire VMR_L4D3_AS_L4D3n3_wr_en;
wire [10:0] AS_L4D3n3_MC_L1L2_L4D3_read_add;
wire [35:0] AS_L4D3n3_MC_L1L2_L4D3;
AllStubs  AS_L4D3n3(
.data_in(VMR_L4D3_AS_L4D3n3),
.enable(VMR_L4D3_AS_L4D3n3_wr_en),
.read_add_MC(AS_L4D3n3_MC_L1L2_L4D3_read_add),
.data_out_MC(AS_L4D3n3_MC_L1L2_L4D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D4PHI1Z1_CM_L1L2_L4D4PHI1Z1;
wire ME_L1L2_L4D4PHI1Z1_CM_L1L2_L4D4PHI1Z1_wr_en;
wire [5:0] CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI1Z1(
.data_in(ME_L1L2_L4D4PHI1Z1_CM_L1L2_L4D4PHI1Z1),
.enable(ME_L1L2_L4D4PHI1Z1_CM_L1L2_L4D4PHI1Z1_wr_en),
.number_out(CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D4PHI1Z2_CM_L1L2_L4D4PHI1Z2;
wire ME_L1L2_L4D4PHI1Z2_CM_L1L2_L4D4PHI1Z2_wr_en;
wire [5:0] CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI1Z2(
.data_in(ME_L1L2_L4D4PHI1Z2_CM_L1L2_L4D4PHI1Z2),
.enable(ME_L1L2_L4D4PHI1Z2_CM_L1L2_L4D4PHI1Z2_wr_en),
.number_out(CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D4PHI2Z1_CM_L1L2_L4D4PHI2Z1;
wire ME_L1L2_L4D4PHI2Z1_CM_L1L2_L4D4PHI2Z1_wr_en;
wire [5:0] CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI2Z1(
.data_in(ME_L1L2_L4D4PHI2Z1_CM_L1L2_L4D4PHI2Z1),
.enable(ME_L1L2_L4D4PHI2Z1_CM_L1L2_L4D4PHI2Z1_wr_en),
.number_out(CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D4PHI2Z2_CM_L1L2_L4D4PHI2Z2;
wire ME_L1L2_L4D4PHI2Z2_CM_L1L2_L4D4PHI2Z2_wr_en;
wire [5:0] CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI2Z2(
.data_in(ME_L1L2_L4D4PHI2Z2_CM_L1L2_L4D4PHI2Z2),
.enable(ME_L1L2_L4D4PHI2Z2_CM_L1L2_L4D4PHI2Z2_wr_en),
.number_out(CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D4PHI3Z1_CM_L1L2_L4D4PHI3Z1;
wire ME_L1L2_L4D4PHI3Z1_CM_L1L2_L4D4PHI3Z1_wr_en;
wire [5:0] CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI3Z1(
.data_in(ME_L1L2_L4D4PHI3Z1_CM_L1L2_L4D4PHI3Z1),
.enable(ME_L1L2_L4D4PHI3Z1_CM_L1L2_L4D4PHI3Z1_wr_en),
.number_out(CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D4PHI3Z2_CM_L1L2_L4D4PHI3Z2;
wire ME_L1L2_L4D4PHI3Z2_CM_L1L2_L4D4PHI3Z2_wr_en;
wire [5:0] CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI3Z2(
.data_in(ME_L1L2_L4D4PHI3Z2_CM_L1L2_L4D4PHI3Z2),
.enable(ME_L1L2_L4D4PHI3Z2_CM_L1L2_L4D4PHI3Z2_wr_en),
.number_out(CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D4PHI4Z1_CM_L1L2_L4D4PHI4Z1;
wire ME_L1L2_L4D4PHI4Z1_CM_L1L2_L4D4PHI4Z1_wr_en;
wire [5:0] CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI4Z1(
.data_in(ME_L1L2_L4D4PHI4Z1_CM_L1L2_L4D4PHI4Z1),
.enable(ME_L1L2_L4D4PHI4Z1_CM_L1L2_L4D4PHI4Z1_wr_en),
.number_out(CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L4D4PHI4Z2_CM_L1L2_L4D4PHI4Z2;
wire ME_L1L2_L4D4PHI4Z2_CM_L1L2_L4D4PHI4Z2_wr_en;
wire [5:0] CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI4Z2(
.data_in(ME_L1L2_L4D4PHI4Z2_CM_L1L2_L4D4PHI4Z2),
.enable(ME_L1L2_L4D4PHI4Z2_CM_L1L2_L4D4PHI4Z2_wr_en),
.number_out(CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L4D4_L1L2_AP_L1L2_L4D4;
wire PR_L4D4_L1L2_AP_L1L2_L4D4_wr_en;
wire [8:0] AP_L1L2_L4D4_MC_L1L2_L4D4_read_add;
wire [55:0] AP_L1L2_L4D4_MC_L1L2_L4D4;
AllProj #(1'b0) AP_L1L2_L4D4(
.data_in(PR_L4D4_L1L2_AP_L1L2_L4D4),
.enable(PR_L4D4_L1L2_AP_L1L2_L4D4_wr_en),
.read_add(AP_L1L2_L4D4_MC_L1L2_L4D4_read_add),
.data_out(AP_L1L2_L4D4_MC_L1L2_L4D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L4D4_AS_L4D4n4;
wire VMR_L4D4_AS_L4D4n4_wr_en;
wire [10:0] AS_L4D4n4_MC_L1L2_L4D4_read_add;
wire [35:0] AS_L4D4n4_MC_L1L2_L4D4;
AllStubs  AS_L4D4n4(
.data_in(VMR_L4D4_AS_L4D4n4),
.enable(VMR_L4D4_AS_L4D4n4_wr_en),
.read_add_MC(AS_L4D4n4_MC_L1L2_L4D4_read_add),
.data_out_MC(AS_L4D4n4_MC_L1L2_L4D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D3PHI1Z1_CM_L1L2_L5D3PHI1Z1;
wire ME_L1L2_L5D3PHI1Z1_CM_L1L2_L5D3PHI1Z1_wr_en;
wire [5:0] CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI1Z1(
.data_in(ME_L1L2_L5D3PHI1Z1_CM_L1L2_L5D3PHI1Z1),
.enable(ME_L1L2_L5D3PHI1Z1_CM_L1L2_L5D3PHI1Z1_wr_en),
.number_out(CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D3PHI1Z2_CM_L1L2_L5D3PHI1Z2;
wire ME_L1L2_L5D3PHI1Z2_CM_L1L2_L5D3PHI1Z2_wr_en;
wire [5:0] CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI1Z2(
.data_in(ME_L1L2_L5D3PHI1Z2_CM_L1L2_L5D3PHI1Z2),
.enable(ME_L1L2_L5D3PHI1Z2_CM_L1L2_L5D3PHI1Z2_wr_en),
.number_out(CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D3PHI2Z1_CM_L1L2_L5D3PHI2Z1;
wire ME_L1L2_L5D3PHI2Z1_CM_L1L2_L5D3PHI2Z1_wr_en;
wire [5:0] CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI2Z1(
.data_in(ME_L1L2_L5D3PHI2Z1_CM_L1L2_L5D3PHI2Z1),
.enable(ME_L1L2_L5D3PHI2Z1_CM_L1L2_L5D3PHI2Z1_wr_en),
.number_out(CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D3PHI2Z2_CM_L1L2_L5D3PHI2Z2;
wire ME_L1L2_L5D3PHI2Z2_CM_L1L2_L5D3PHI2Z2_wr_en;
wire [5:0] CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI2Z2(
.data_in(ME_L1L2_L5D3PHI2Z2_CM_L1L2_L5D3PHI2Z2),
.enable(ME_L1L2_L5D3PHI2Z2_CM_L1L2_L5D3PHI2Z2_wr_en),
.number_out(CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D3PHI3Z1_CM_L1L2_L5D3PHI3Z1;
wire ME_L1L2_L5D3PHI3Z1_CM_L1L2_L5D3PHI3Z1_wr_en;
wire [5:0] CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI3Z1(
.data_in(ME_L1L2_L5D3PHI3Z1_CM_L1L2_L5D3PHI3Z1),
.enable(ME_L1L2_L5D3PHI3Z1_CM_L1L2_L5D3PHI3Z1_wr_en),
.number_out(CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D3PHI3Z2_CM_L1L2_L5D3PHI3Z2;
wire ME_L1L2_L5D3PHI3Z2_CM_L1L2_L5D3PHI3Z2_wr_en;
wire [5:0] CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI3Z2(
.data_in(ME_L1L2_L5D3PHI3Z2_CM_L1L2_L5D3PHI3Z2),
.enable(ME_L1L2_L5D3PHI3Z2_CM_L1L2_L5D3PHI3Z2_wr_en),
.number_out(CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L5D3_L1L2_AP_L1L2_L5D3;
wire PR_L5D3_L1L2_AP_L1L2_L5D3_wr_en;
wire [8:0] AP_L1L2_L5D3_MC_L1L2_L5D3_read_add;
wire [55:0] AP_L1L2_L5D3_MC_L1L2_L5D3;
AllProj #(1'b0) AP_L1L2_L5D3(
.data_in(PR_L5D3_L1L2_AP_L1L2_L5D3),
.enable(PR_L5D3_L1L2_AP_L1L2_L5D3_wr_en),
.read_add(AP_L1L2_L5D3_MC_L1L2_L5D3_read_add),
.data_out(AP_L1L2_L5D3_MC_L1L2_L5D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L5D3_AS_L5D3n4;
wire VMR_L5D3_AS_L5D3n4_wr_en;
wire [10:0] AS_L5D3n4_MC_L1L2_L5D3_read_add;
wire [35:0] AS_L5D3n4_MC_L1L2_L5D3;
AllStubs  AS_L5D3n4(
.data_in(VMR_L5D3_AS_L5D3n4),
.enable(VMR_L5D3_AS_L5D3n4_wr_en),
.read_add_MC(AS_L5D3n4_MC_L1L2_L5D3_read_add),
.data_out_MC(AS_L5D3n4_MC_L1L2_L5D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D4PHI1Z1_CM_L1L2_L5D4PHI1Z1;
wire ME_L1L2_L5D4PHI1Z1_CM_L1L2_L5D4PHI1Z1_wr_en;
wire [5:0] CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI1Z1(
.data_in(ME_L1L2_L5D4PHI1Z1_CM_L1L2_L5D4PHI1Z1),
.enable(ME_L1L2_L5D4PHI1Z1_CM_L1L2_L5D4PHI1Z1_wr_en),
.number_out(CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D4PHI1Z2_CM_L1L2_L5D4PHI1Z2;
wire ME_L1L2_L5D4PHI1Z2_CM_L1L2_L5D4PHI1Z2_wr_en;
wire [5:0] CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI1Z2(
.data_in(ME_L1L2_L5D4PHI1Z2_CM_L1L2_L5D4PHI1Z2),
.enable(ME_L1L2_L5D4PHI1Z2_CM_L1L2_L5D4PHI1Z2_wr_en),
.number_out(CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D4PHI2Z1_CM_L1L2_L5D4PHI2Z1;
wire ME_L1L2_L5D4PHI2Z1_CM_L1L2_L5D4PHI2Z1_wr_en;
wire [5:0] CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI2Z1(
.data_in(ME_L1L2_L5D4PHI2Z1_CM_L1L2_L5D4PHI2Z1),
.enable(ME_L1L2_L5D4PHI2Z1_CM_L1L2_L5D4PHI2Z1_wr_en),
.number_out(CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D4PHI2Z2_CM_L1L2_L5D4PHI2Z2;
wire ME_L1L2_L5D4PHI2Z2_CM_L1L2_L5D4PHI2Z2_wr_en;
wire [5:0] CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI2Z2(
.data_in(ME_L1L2_L5D4PHI2Z2_CM_L1L2_L5D4PHI2Z2),
.enable(ME_L1L2_L5D4PHI2Z2_CM_L1L2_L5D4PHI2Z2_wr_en),
.number_out(CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D4PHI3Z1_CM_L1L2_L5D4PHI3Z1;
wire ME_L1L2_L5D4PHI3Z1_CM_L1L2_L5D4PHI3Z1_wr_en;
wire [5:0] CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI3Z1(
.data_in(ME_L1L2_L5D4PHI3Z1_CM_L1L2_L5D4PHI3Z1),
.enable(ME_L1L2_L5D4PHI3Z1_CM_L1L2_L5D4PHI3Z1_wr_en),
.number_out(CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L5D4PHI3Z2_CM_L1L2_L5D4PHI3Z2;
wire ME_L1L2_L5D4PHI3Z2_CM_L1L2_L5D4PHI3Z2_wr_en;
wire [5:0] CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI3Z2(
.data_in(ME_L1L2_L5D4PHI3Z2_CM_L1L2_L5D4PHI3Z2),
.enable(ME_L1L2_L5D4PHI3Z2_CM_L1L2_L5D4PHI3Z2_wr_en),
.number_out(CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L5D4_L1L2_AP_L1L2_L5D4;
wire PR_L5D4_L1L2_AP_L1L2_L5D4_wr_en;
wire [8:0] AP_L1L2_L5D4_MC_L1L2_L5D4_read_add;
wire [55:0] AP_L1L2_L5D4_MC_L1L2_L5D4;
AllProj #(1'b0) AP_L1L2_L5D4(
.data_in(PR_L5D4_L1L2_AP_L1L2_L5D4),
.enable(PR_L5D4_L1L2_AP_L1L2_L5D4_wr_en),
.read_add(AP_L1L2_L5D4_MC_L1L2_L5D4_read_add),
.data_out(AP_L1L2_L5D4_MC_L1L2_L5D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L5D4_AS_L5D4n3;
wire VMR_L5D4_AS_L5D4n3_wr_en;
wire [10:0] AS_L5D4n3_MC_L1L2_L5D4_read_add;
wire [35:0] AS_L5D4n3_MC_L1L2_L5D4;
AllStubs  AS_L5D4n3(
.data_in(VMR_L5D4_AS_L5D4n3),
.enable(VMR_L5D4_AS_L5D4n3_wr_en),
.read_add_MC(AS_L5D4n3_MC_L1L2_L5D4_read_add),
.data_out_MC(AS_L5D4n3_MC_L1L2_L5D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D3PHI1Z1_CM_L1L2_L6D3PHI1Z1;
wire ME_L1L2_L6D3PHI1Z1_CM_L1L2_L6D3PHI1Z1_wr_en;
wire [5:0] CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI1Z1(
.data_in(ME_L1L2_L6D3PHI1Z1_CM_L1L2_L6D3PHI1Z1),
.enable(ME_L1L2_L6D3PHI1Z1_CM_L1L2_L6D3PHI1Z1_wr_en),
.number_out(CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D3PHI1Z2_CM_L1L2_L6D3PHI1Z2;
wire ME_L1L2_L6D3PHI1Z2_CM_L1L2_L6D3PHI1Z2_wr_en;
wire [5:0] CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI1Z2(
.data_in(ME_L1L2_L6D3PHI1Z2_CM_L1L2_L6D3PHI1Z2),
.enable(ME_L1L2_L6D3PHI1Z2_CM_L1L2_L6D3PHI1Z2_wr_en),
.number_out(CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D3PHI2Z1_CM_L1L2_L6D3PHI2Z1;
wire ME_L1L2_L6D3PHI2Z1_CM_L1L2_L6D3PHI2Z1_wr_en;
wire [5:0] CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI2Z1(
.data_in(ME_L1L2_L6D3PHI2Z1_CM_L1L2_L6D3PHI2Z1),
.enable(ME_L1L2_L6D3PHI2Z1_CM_L1L2_L6D3PHI2Z1_wr_en),
.number_out(CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D3PHI2Z2_CM_L1L2_L6D3PHI2Z2;
wire ME_L1L2_L6D3PHI2Z2_CM_L1L2_L6D3PHI2Z2_wr_en;
wire [5:0] CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI2Z2(
.data_in(ME_L1L2_L6D3PHI2Z2_CM_L1L2_L6D3PHI2Z2),
.enable(ME_L1L2_L6D3PHI2Z2_CM_L1L2_L6D3PHI2Z2_wr_en),
.number_out(CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D3PHI3Z1_CM_L1L2_L6D3PHI3Z1;
wire ME_L1L2_L6D3PHI3Z1_CM_L1L2_L6D3PHI3Z1_wr_en;
wire [5:0] CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI3Z1(
.data_in(ME_L1L2_L6D3PHI3Z1_CM_L1L2_L6D3PHI3Z1),
.enable(ME_L1L2_L6D3PHI3Z1_CM_L1L2_L6D3PHI3Z1_wr_en),
.number_out(CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D3PHI3Z2_CM_L1L2_L6D3PHI3Z2;
wire ME_L1L2_L6D3PHI3Z2_CM_L1L2_L6D3PHI3Z2_wr_en;
wire [5:0] CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI3Z2(
.data_in(ME_L1L2_L6D3PHI3Z2_CM_L1L2_L6D3PHI3Z2),
.enable(ME_L1L2_L6D3PHI3Z2_CM_L1L2_L6D3PHI3Z2_wr_en),
.number_out(CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D3PHI4Z1_CM_L1L2_L6D3PHI4Z1;
wire ME_L1L2_L6D3PHI4Z1_CM_L1L2_L6D3PHI4Z1_wr_en;
wire [5:0] CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI4Z1(
.data_in(ME_L1L2_L6D3PHI4Z1_CM_L1L2_L6D3PHI4Z1),
.enable(ME_L1L2_L6D3PHI4Z1_CM_L1L2_L6D3PHI4Z1_wr_en),
.number_out(CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D3PHI4Z2_CM_L1L2_L6D3PHI4Z2;
wire ME_L1L2_L6D3PHI4Z2_CM_L1L2_L6D3PHI4Z2_wr_en;
wire [5:0] CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI4Z2(
.data_in(ME_L1L2_L6D3PHI4Z2_CM_L1L2_L6D3PHI4Z2),
.enable(ME_L1L2_L6D3PHI4Z2_CM_L1L2_L6D3PHI4Z2_wr_en),
.number_out(CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L6D3_L1L2_AP_L1L2_L6D3;
wire PR_L6D3_L1L2_AP_L1L2_L6D3_wr_en;
wire [8:0] AP_L1L2_L6D3_MC_L1L2_L6D3_read_add;
wire [55:0] AP_L1L2_L6D3_MC_L1L2_L6D3;
AllProj #(1'b0) AP_L1L2_L6D3(
.data_in(PR_L6D3_L1L2_AP_L1L2_L6D3),
.enable(PR_L6D3_L1L2_AP_L1L2_L6D3_wr_en),
.read_add(AP_L1L2_L6D3_MC_L1L2_L6D3_read_add),
.data_out(AP_L1L2_L6D3_MC_L1L2_L6D3),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L6D3_AS_L6D3n3;
wire VMR_L6D3_AS_L6D3n3_wr_en;
wire [10:0] AS_L6D3n3_MC_L1L2_L6D3_read_add;
wire [35:0] AS_L6D3n3_MC_L1L2_L6D3;
AllStubs  AS_L6D3n3(
.data_in(VMR_L6D3_AS_L6D3n3),
.enable(VMR_L6D3_AS_L6D3n3_wr_en),
.read_add_MC(AS_L6D3n3_MC_L1L2_L6D3_read_add),
.data_out_MC(AS_L6D3n3_MC_L1L2_L6D3),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D4PHI1Z1_CM_L1L2_L6D4PHI1Z1;
wire ME_L1L2_L6D4PHI1Z1_CM_L1L2_L6D4PHI1Z1_wr_en;
wire [5:0] CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI1Z1(
.data_in(ME_L1L2_L6D4PHI1Z1_CM_L1L2_L6D4PHI1Z1),
.enable(ME_L1L2_L6D4PHI1Z1_CM_L1L2_L6D4PHI1Z1_wr_en),
.number_out(CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D4PHI1Z2_CM_L1L2_L6D4PHI1Z2;
wire ME_L1L2_L6D4PHI1Z2_CM_L1L2_L6D4PHI1Z2_wr_en;
wire [5:0] CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI1Z2(
.data_in(ME_L1L2_L6D4PHI1Z2_CM_L1L2_L6D4PHI1Z2),
.enable(ME_L1L2_L6D4PHI1Z2_CM_L1L2_L6D4PHI1Z2_wr_en),
.number_out(CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D4PHI2Z1_CM_L1L2_L6D4PHI2Z1;
wire ME_L1L2_L6D4PHI2Z1_CM_L1L2_L6D4PHI2Z1_wr_en;
wire [5:0] CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI2Z1(
.data_in(ME_L1L2_L6D4PHI2Z1_CM_L1L2_L6D4PHI2Z1),
.enable(ME_L1L2_L6D4PHI2Z1_CM_L1L2_L6D4PHI2Z1_wr_en),
.number_out(CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D4PHI2Z2_CM_L1L2_L6D4PHI2Z2;
wire ME_L1L2_L6D4PHI2Z2_CM_L1L2_L6D4PHI2Z2_wr_en;
wire [5:0] CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI2Z2(
.data_in(ME_L1L2_L6D4PHI2Z2_CM_L1L2_L6D4PHI2Z2),
.enable(ME_L1L2_L6D4PHI2Z2_CM_L1L2_L6D4PHI2Z2_wr_en),
.number_out(CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D4PHI3Z1_CM_L1L2_L6D4PHI3Z1;
wire ME_L1L2_L6D4PHI3Z1_CM_L1L2_L6D4PHI3Z1_wr_en;
wire [5:0] CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI3Z1(
.data_in(ME_L1L2_L6D4PHI3Z1_CM_L1L2_L6D4PHI3Z1),
.enable(ME_L1L2_L6D4PHI3Z1_CM_L1L2_L6D4PHI3Z1_wr_en),
.number_out(CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D4PHI3Z2_CM_L1L2_L6D4PHI3Z2;
wire ME_L1L2_L6D4PHI3Z2_CM_L1L2_L6D4PHI3Z2_wr_en;
wire [5:0] CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI3Z2(
.data_in(ME_L1L2_L6D4PHI3Z2_CM_L1L2_L6D4PHI3Z2),
.enable(ME_L1L2_L6D4PHI3Z2_CM_L1L2_L6D4PHI3Z2_wr_en),
.number_out(CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D4PHI4Z1_CM_L1L2_L6D4PHI4Z1;
wire ME_L1L2_L6D4PHI4Z1_CM_L1L2_L6D4PHI4Z1_wr_en;
wire [5:0] CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI4Z1(
.data_in(ME_L1L2_L6D4PHI4Z1_CM_L1L2_L6D4PHI4Z1),
.enable(ME_L1L2_L6D4PHI4Z1_CM_L1L2_L6D4PHI4Z1_wr_en),
.number_out(CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [11:0] ME_L1L2_L6D4PHI4Z2_CM_L1L2_L6D4PHI4Z2;
wire ME_L1L2_L6D4PHI4Z2_CM_L1L2_L6D4PHI4Z2_wr_en;
wire [5:0] CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI4Z2(
.data_in(ME_L1L2_L6D4PHI4Z2_CM_L1L2_L6D4PHI4Z2),
.enable(ME_L1L2_L6D4PHI4Z2_CM_L1L2_L6D4PHI4Z2_wr_en),
.number_out(CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4),
.start(start8_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] PR_L6D4_L1L2_AP_L1L2_L6D4;
wire PR_L6D4_L1L2_AP_L1L2_L6D4_wr_en;
wire [8:0] AP_L1L2_L6D4_MC_L1L2_L6D4_read_add;
wire [55:0] AP_L1L2_L6D4_MC_L1L2_L6D4;
AllProj #(1'b0) AP_L1L2_L6D4(
.data_in(PR_L6D4_L1L2_AP_L1L2_L6D4),
.enable(PR_L6D4_L1L2_AP_L1L2_L6D4_wr_en),
.read_add(AP_L1L2_L6D4_MC_L1L2_L6D4_read_add),
.data_out(AP_L1L2_L6D4_MC_L1L2_L6D4),
.start(start7_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] VMR_L6D4_AS_L6D4n4;
wire VMR_L6D4_AS_L6D4n4_wr_en;
wire [10:0] AS_L6D4n4_MC_L1L2_L6D4_read_add;
wire [35:0] AS_L6D4n4_MC_L1L2_L6D4;
AllStubs  AS_L6D4n4(
.data_in(VMR_L6D4_AS_L6D4n4),
.enable(VMR_L6D4_AS_L6D4n4_wr_en),
.read_add_MC(AS_L6D4n4_MC_L1L2_L6D4_read_add),
.data_out_MC(AS_L6D4n4_MC_L1L2_L6D4),
.start(start3_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus;
wire MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus_wr_en;
wire [5:0] FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus_number;
wire [9:0] FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus_read_add;
wire [35:0] FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus;
FullMatch #(128) FM_L3L4_L1D3_ToMinus(
.data_in(MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus),
.enable(MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus_wr_en),
.number_out(FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus_number),
.read_add(FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus_read_add),
.data_out(FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus;
wire MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus_wr_en;
wire [5:0] FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus_number;
wire [9:0] FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus_read_add;
wire [35:0] FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus;
FullMatch #(128) FM_L3L4_L1D4_ToMinus(
.data_in(MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus),
.enable(MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus_wr_en),
.number_out(FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus_number),
.read_add(FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus_read_add),
.data_out(FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus;
wire MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus_wr_en;
wire [5:0] FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus_number;
wire [9:0] FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus_read_add;
wire [35:0] FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus;
FullMatch #(128) FM_L3L4_L2D3_ToMinus(
.data_in(MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus),
.enable(MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus_wr_en),
.number_out(FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus_number),
.read_add(FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus_read_add),
.data_out(FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus;
wire MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus_wr_en;
wire [5:0] FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus_number;
wire [9:0] FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus_read_add;
wire [35:0] FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus;
FullMatch #(128) FM_L3L4_L2D4_ToMinus(
.data_in(MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus),
.enable(MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus_wr_en),
.number_out(FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus_number),
.read_add(FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus_read_add),
.data_out(FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus;
wire MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus_wr_en;
wire [5:0] FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus_number;
wire [9:0] FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus_read_add;
wire [35:0] FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus;
FullMatch #(128) FM_L3L4_L5D3_ToMinus(
.data_in(MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus),
.enable(MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus_wr_en),
.number_out(FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus_number),
.read_add(FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus_read_add),
.data_out(FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus;
wire MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus_wr_en;
wire [5:0] FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus_number;
wire [9:0] FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus_read_add;
wire [35:0] FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus;
FullMatch #(128) FM_L3L4_L5D4_ToMinus(
.data_in(MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus),
.enable(MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus_wr_en),
.number_out(FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus_number),
.read_add(FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus_read_add),
.data_out(FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus;
wire MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus_wr_en;
wire [5:0] FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus_number;
wire [9:0] FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus_read_add;
wire [35:0] FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus;
FullMatch #(128) FM_L3L4_L6D3_ToMinus(
.data_in(MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus),
.enable(MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus_wr_en),
.number_out(FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus_number),
.read_add(FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus_read_add),
.data_out(FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus;
wire MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus_wr_en;
wire [5:0] FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus_number;
wire [9:0] FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus_read_add;
wire [35:0] FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus;
FullMatch #(128) FM_L3L4_L6D4_ToMinus(
.data_in(MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus),
.enable(MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus_wr_en),
.number_out(FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus_number),
.read_add(FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus_read_add),
.data_out(FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus;
wire MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus_wr_en;
wire [5:0] FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus_number;
wire [9:0] FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus_read_add;
wire [35:0] FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus;
FullMatch #(128) FM_L5L6_L1D3_ToMinus(
.data_in(MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus),
.enable(MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus_wr_en),
.number_out(FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus_number),
.read_add(FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus_read_add),
.data_out(FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus;
wire MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus_wr_en;
wire [5:0] FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus_number;
wire [9:0] FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus_read_add;
wire [35:0] FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus;
FullMatch #(128) FM_L5L6_L1D4_ToMinus(
.data_in(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus),
.enable(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus_wr_en),
.number_out(FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus_number),
.read_add(FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus_read_add),
.data_out(FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus;
wire MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus_wr_en;
wire [5:0] FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus_number;
wire [9:0] FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus_read_add;
wire [35:0] FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus;
FullMatch #(128) FM_L5L6_L2D3_ToMinus(
.data_in(MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus),
.enable(MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus_wr_en),
.number_out(FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus_number),
.read_add(FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus_read_add),
.data_out(FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus;
wire MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus_wr_en;
wire [5:0] FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus_number;
wire [9:0] FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus_read_add;
wire [35:0] FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus;
FullMatch #(128) FM_L5L6_L2D4_ToMinus(
.data_in(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus),
.enable(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus_wr_en),
.number_out(FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus_number),
.read_add(FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus_read_add),
.data_out(FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus;
wire MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus_wr_en;
wire [5:0] FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus_number;
wire [9:0] FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus_read_add;
wire [35:0] FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus;
FullMatch #(128) FM_L5L6_L3D3_ToMinus(
.data_in(MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus),
.enable(MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus_wr_en),
.number_out(FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus_number),
.read_add(FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus_read_add),
.data_out(FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus;
wire MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus_wr_en;
wire [5:0] FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus_number;
wire [9:0] FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus_read_add;
wire [35:0] FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus;
FullMatch #(128) FM_L5L6_L3D4_ToMinus(
.data_in(MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus),
.enable(MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus_wr_en),
.number_out(FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus_number),
.read_add(FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus_read_add),
.data_out(FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus;
wire MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus_wr_en;
wire [5:0] FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus_number;
wire [9:0] FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus_read_add;
wire [35:0] FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus;
FullMatch #(128) FM_L5L6_L4D3_ToMinus(
.data_in(MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus),
.enable(MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus_wr_en),
.number_out(FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus_number),
.read_add(FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus_read_add),
.data_out(FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus;
wire MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus_wr_en;
wire [5:0] FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus_number;
wire [9:0] FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus_read_add;
wire [35:0] FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus;
FullMatch #(128) FM_L5L6_L4D4_ToMinus(
.data_in(MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus),
.enable(MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus_wr_en),
.number_out(FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus_number),
.read_add(FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus_read_add),
.data_out(FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus;
wire MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus_wr_en;
wire [5:0] FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus_number;
wire [9:0] FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus_read_add;
wire [35:0] FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus;
FullMatch #(128) FM_L1L2_L3D3_ToMinus(
.data_in(MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus),
.enable(MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus_wr_en),
.number_out(FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus_number),
.read_add(FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus_read_add),
.data_out(FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus;
wire MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus_wr_en;
wire [5:0] FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus_number;
wire [9:0] FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus_read_add;
wire [35:0] FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus;
FullMatch #(128) FM_L1L2_L3D4_ToMinus(
.data_in(MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus),
.enable(MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus_wr_en),
.number_out(FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus_number),
.read_add(FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus_read_add),
.data_out(FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus;
wire MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus_wr_en;
wire [5:0] FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus_number;
wire [9:0] FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus_read_add;
wire [35:0] FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus;
FullMatch #(128) FM_L1L2_L4D3_ToMinus(
.data_in(MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus),
.enable(MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus_wr_en),
.number_out(FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus_number),
.read_add(FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus_read_add),
.data_out(FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus;
wire MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus_wr_en;
wire [5:0] FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus_number;
wire [9:0] FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus_read_add;
wire [35:0] FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus;
FullMatch #(128) FM_L1L2_L4D4_ToMinus(
.data_in(MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus),
.enable(MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus_wr_en),
.number_out(FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus_number),
.read_add(FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus_read_add),
.data_out(FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus;
wire MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus_wr_en;
wire [5:0] FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus_number;
wire [9:0] FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus_read_add;
wire [35:0] FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus;
FullMatch #(128) FM_L1L2_L5D3_ToMinus(
.data_in(MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus),
.enable(MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus_wr_en),
.number_out(FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus_number),
.read_add(FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus_read_add),
.data_out(FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus;
wire MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus_wr_en;
wire [5:0] FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus_number;
wire [9:0] FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus_read_add;
wire [35:0] FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus;
FullMatch #(128) FM_L1L2_L5D4_ToMinus(
.data_in(MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus),
.enable(MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus_wr_en),
.number_out(FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus_number),
.read_add(FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus_read_add),
.data_out(FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus;
wire MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus_wr_en;
wire [5:0] FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus_number;
wire [9:0] FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus_read_add;
wire [35:0] FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus;
FullMatch #(128) FM_L1L2_L6D3_ToMinus(
.data_in(MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus),
.enable(MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus_wr_en),
.number_out(FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus_number),
.read_add(FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus_read_add),
.data_out(FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus;
wire MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus_wr_en;
wire [5:0] FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus_number;
wire [9:0] FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus_read_add;
wire [35:0] FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus;
FullMatch #(128) FM_L1L2_L6D4_ToMinus(
.data_in(MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus),
.enable(MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus_wr_en),
.number_out(FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus_number),
.read_add(FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus_read_add),
.data_out(FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus;
wire MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus_wr_en;
wire [5:0] FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus_number;
wire [9:0] FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus_read_add;
wire [35:0] FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus;
FullMatch #(128) FM_L3L4_L1D3_ToPlus(
.data_in(MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus),
.enable(MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus_wr_en),
.number_out(FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus_number),
.read_add(FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus_read_add),
.data_out(FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus;
wire MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus_wr_en;
wire [5:0] FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus_number;
wire [9:0] FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus_read_add;
wire [35:0] FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus;
FullMatch #(128) FM_L3L4_L1D4_ToPlus(
.data_in(MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus),
.enable(MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus_wr_en),
.number_out(FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus_number),
.read_add(FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus_read_add),
.data_out(FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus;
wire MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus_wr_en;
wire [5:0] FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus_number;
wire [9:0] FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus_read_add;
wire [35:0] FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus;
FullMatch #(128) FM_L3L4_L2D3_ToPlus(
.data_in(MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus),
.enable(MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus_wr_en),
.number_out(FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus_number),
.read_add(FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus_read_add),
.data_out(FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus;
wire MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus_wr_en;
wire [5:0] FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus_number;
wire [9:0] FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus_read_add;
wire [35:0] FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus;
FullMatch #(128) FM_L3L4_L2D4_ToPlus(
.data_in(MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus),
.enable(MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus_wr_en),
.number_out(FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus_number),
.read_add(FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus_read_add),
.data_out(FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus;
wire MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus_wr_en;
wire [5:0] FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus_number;
wire [9:0] FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus_read_add;
wire [35:0] FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus;
FullMatch #(128) FM_L3L4_L5D3_ToPlus(
.data_in(MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus),
.enable(MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus_wr_en),
.number_out(FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus_number),
.read_add(FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus_read_add),
.data_out(FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus;
wire MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus_wr_en;
wire [5:0] FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus_number;
wire [9:0] FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus_read_add;
wire [35:0] FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus;
FullMatch #(128) FM_L3L4_L5D4_ToPlus(
.data_in(MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus),
.enable(MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus_wr_en),
.number_out(FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus_number),
.read_add(FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus_read_add),
.data_out(FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus;
wire MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus_wr_en;
wire [5:0] FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus_number;
wire [9:0] FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus_read_add;
wire [35:0] FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus;
FullMatch #(128) FM_L3L4_L6D3_ToPlus(
.data_in(MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus),
.enable(MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus_wr_en),
.number_out(FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus_number),
.read_add(FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus_read_add),
.data_out(FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus;
wire MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus_wr_en;
wire [5:0] FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus_number;
wire [9:0] FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus_read_add;
wire [35:0] FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus;
FullMatch #(128) FM_L3L4_L6D4_ToPlus(
.data_in(MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus),
.enable(MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus_wr_en),
.number_out(FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus_number),
.read_add(FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus_read_add),
.data_out(FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus;
wire MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus_wr_en;
wire [5:0] FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus_number;
wire [9:0] FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus_read_add;
wire [35:0] FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus;
FullMatch #(128) FM_L5L6_L1D3_ToPlus(
.data_in(MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus),
.enable(MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus_wr_en),
.number_out(FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus_number),
.read_add(FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus_read_add),
.data_out(FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus;
wire MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus_wr_en;
wire [5:0] FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus_number;
wire [9:0] FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus_read_add;
wire [35:0] FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus;
FullMatch #(128) FM_L5L6_L1D4_ToPlus(
.data_in(MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus),
.enable(MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus_wr_en),
.number_out(FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus_number),
.read_add(FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus_read_add),
.data_out(FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus;
wire MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus_wr_en;
wire [5:0] FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus_number;
wire [9:0] FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus_read_add;
wire [35:0] FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus;
FullMatch #(128) FM_L5L6_L2D3_ToPlus(
.data_in(MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus),
.enable(MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus_wr_en),
.number_out(FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus_number),
.read_add(FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus_read_add),
.data_out(FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus;
wire MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus_wr_en;
wire [5:0] FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus_number;
wire [9:0] FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus_read_add;
wire [35:0] FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus;
FullMatch #(128) FM_L5L6_L2D4_ToPlus(
.data_in(MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus),
.enable(MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus_wr_en),
.number_out(FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus_number),
.read_add(FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus_read_add),
.data_out(FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus;
wire MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus_wr_en;
wire [5:0] FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus_number;
wire [9:0] FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus_read_add;
wire [35:0] FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus;
FullMatch #(128) FM_L5L6_L3D3_ToPlus(
.data_in(MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus),
.enable(MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus_wr_en),
.number_out(FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus_number),
.read_add(FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus_read_add),
.data_out(FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus;
wire MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus_wr_en;
wire [5:0] FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus_number;
wire [9:0] FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus_read_add;
wire [35:0] FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus;
FullMatch #(128) FM_L5L6_L3D4_ToPlus(
.data_in(MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus),
.enable(MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus_wr_en),
.number_out(FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus_number),
.read_add(FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus_read_add),
.data_out(FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus;
wire MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus_wr_en;
wire [5:0] FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus_number;
wire [9:0] FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus_read_add;
wire [35:0] FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus;
FullMatch #(128) FM_L5L6_L4D3_ToPlus(
.data_in(MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus),
.enable(MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus_wr_en),
.number_out(FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus_number),
.read_add(FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus_read_add),
.data_out(FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus;
wire MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus_wr_en;
wire [5:0] FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus_number;
wire [9:0] FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus_read_add;
wire [35:0] FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus;
FullMatch #(128) FM_L5L6_L4D4_ToPlus(
.data_in(MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus),
.enable(MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus_wr_en),
.number_out(FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus_number),
.read_add(FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus_read_add),
.data_out(FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus;
wire MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus_wr_en;
wire [5:0] FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus_number;
wire [9:0] FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus_read_add;
wire [35:0] FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus;
FullMatch #(128) FM_L1L2_L3D3_ToPlus(
.data_in(MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus),
.enable(MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus_wr_en),
.number_out(FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus_number),
.read_add(FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus_read_add),
.data_out(FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus;
wire MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus_wr_en;
wire [5:0] FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus_number;
wire [9:0] FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus_read_add;
wire [35:0] FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus;
FullMatch #(128) FM_L1L2_L3D4_ToPlus(
.data_in(MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus),
.enable(MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus_wr_en),
.number_out(FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus_number),
.read_add(FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus_read_add),
.data_out(FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus;
wire MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus_wr_en;
wire [5:0] FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus_number;
wire [9:0] FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus_read_add;
wire [35:0] FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus;
FullMatch #(128) FM_L1L2_L4D3_ToPlus(
.data_in(MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus),
.enable(MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus_wr_en),
.number_out(FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus_number),
.read_add(FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus_read_add),
.data_out(FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus;
wire MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus_wr_en;
wire [5:0] FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus_number;
wire [9:0] FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus_read_add;
wire [35:0] FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus;
FullMatch #(128) FM_L1L2_L4D4_ToPlus(
.data_in(MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus),
.enable(MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus_wr_en),
.number_out(FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus_number),
.read_add(FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus_read_add),
.data_out(FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus;
wire MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus_wr_en;
wire [5:0] FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus_number;
wire [9:0] FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus_read_add;
wire [35:0] FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus;
FullMatch #(128) FM_L1L2_L5D3_ToPlus(
.data_in(MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus),
.enable(MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus_wr_en),
.number_out(FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus_number),
.read_add(FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus_read_add),
.data_out(FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus;
wire MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus_wr_en;
wire [5:0] FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus_number;
wire [9:0] FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus_read_add;
wire [35:0] FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus;
FullMatch #(128) FM_L1L2_L5D4_ToPlus(
.data_in(MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus),
.enable(MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus_wr_en),
.number_out(FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus_number),
.read_add(FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus_read_add),
.data_out(FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus;
wire MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus_wr_en;
wire [5:0] FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus_number;
wire [9:0] FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus_read_add;
wire [35:0] FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus;
FullMatch #(128) FM_L1L2_L6D3_ToPlus(
.data_in(MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus),
.enable(MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus_wr_en),
.number_out(FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus_number),
.read_add(FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus_read_add),
.data_out(FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus;
wire MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus_wr_en;
wire [5:0] FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus_number;
wire [9:0] FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus_read_add;
wire [35:0] FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus;
FullMatch #(128) FM_L1L2_L6D4_ToPlus(
.data_in(MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus),
.enable(MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus_wr_en),
.number_out(FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus_number),
.read_add(FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus_read_add),
.data_out(FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus),
.read_en(1'b1),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L3D3_FM_L1L2_L3D3;
wire MC_L1L2_L3D3_FM_L1L2_L3D3_wr_en;
wire [5:0] FM_L1L2_L3D3_FT_L1L2_number;
wire [9:0] FM_L1L2_L3D3_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L3D3_FT_L1L2;
wire FM_L1L2_L3D3_FT_L1L2_read_en;
FullMatch  FM_L1L2_L3D3(
.data_in(MC_L1L2_L3D3_FM_L1L2_L3D3),
.enable(MC_L1L2_L3D3_FM_L1L2_L3D3_wr_en),
.number_out(FM_L1L2_L3D3_FT_L1L2_number),
.read_add(FM_L1L2_L3D3_FT_L1L2_read_add),
.data_out(FM_L1L2_L3D3_FT_L1L2),
.read_en(FM_L1L2_L3D3_FT_L1L2_read_en),
.start(start9_0),
.done(done8_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L3D4_FM_L1L2_L3D4;
wire MC_L1L2_L3D4_FM_L1L2_L3D4_wr_en;
wire [5:0] FM_L1L2_L3D4_FT_L1L2_number;
wire [9:0] FM_L1L2_L3D4_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L3D4_FT_L1L2;
wire FM_L1L2_L3D4_FT_L1L2_read_en;
FullMatch  FM_L1L2_L3D4(
.data_in(MC_L1L2_L3D4_FM_L1L2_L3D4),
.enable(MC_L1L2_L3D4_FM_L1L2_L3D4_wr_en),
.number_out(FM_L1L2_L3D4_FT_L1L2_number),
.read_add(FM_L1L2_L3D4_FT_L1L2_read_add),
.data_out(FM_L1L2_L3D4_FT_L1L2),
.read_en(FM_L1L2_L3D4_FT_L1L2_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L4D3_FM_L1L2_L4D3;
wire MC_L1L2_L4D3_FM_L1L2_L4D3_wr_en;
wire [5:0] FM_L1L2_L4D3_FT_L1L2_number;
wire [9:0] FM_L1L2_L4D3_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L4D3_FT_L1L2;
wire FM_L1L2_L4D3_FT_L1L2_read_en;
FullMatch  FM_L1L2_L4D3(
.data_in(MC_L1L2_L4D3_FM_L1L2_L4D3),
.enable(MC_L1L2_L4D3_FM_L1L2_L4D3_wr_en),
.number_out(FM_L1L2_L4D3_FT_L1L2_number),
.read_add(FM_L1L2_L4D3_FT_L1L2_read_add),
.data_out(FM_L1L2_L4D3_FT_L1L2),
.read_en(FM_L1L2_L4D3_FT_L1L2_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L4D4_FM_L1L2_L4D4;
wire MC_L1L2_L4D4_FM_L1L2_L4D4_wr_en;
wire [5:0] FM_L1L2_L4D4_FT_L1L2_number;
wire [9:0] FM_L1L2_L4D4_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L4D4_FT_L1L2;
wire FM_L1L2_L4D4_FT_L1L2_read_en;
FullMatch  FM_L1L2_L4D4(
.data_in(MC_L1L2_L4D4_FM_L1L2_L4D4),
.enable(MC_L1L2_L4D4_FM_L1L2_L4D4_wr_en),
.number_out(FM_L1L2_L4D4_FT_L1L2_number),
.read_add(FM_L1L2_L4D4_FT_L1L2_read_add),
.data_out(FM_L1L2_L4D4_FT_L1L2),
.read_en(FM_L1L2_L4D4_FT_L1L2_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L5D3_FM_L1L2_L5D3;
wire MC_L1L2_L5D3_FM_L1L2_L5D3_wr_en;
wire [5:0] FM_L1L2_L5D3_FT_L1L2_number;
wire [9:0] FM_L1L2_L5D3_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L5D3_FT_L1L2;
wire FM_L1L2_L5D3_FT_L1L2_read_en;
FullMatch  FM_L1L2_L5D3(
.data_in(MC_L1L2_L5D3_FM_L1L2_L5D3),
.enable(MC_L1L2_L5D3_FM_L1L2_L5D3_wr_en),
.number_out(FM_L1L2_L5D3_FT_L1L2_number),
.read_add(FM_L1L2_L5D3_FT_L1L2_read_add),
.data_out(FM_L1L2_L5D3_FT_L1L2),
.read_en(FM_L1L2_L5D3_FT_L1L2_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L5D4_FM_L1L2_L5D4;
wire MC_L1L2_L5D4_FM_L1L2_L5D4_wr_en;
wire [5:0] FM_L1L2_L5D4_FT_L1L2_number;
wire [9:0] FM_L1L2_L5D4_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L5D4_FT_L1L2;
wire FM_L1L2_L5D4_FT_L1L2_read_en;
FullMatch  FM_L1L2_L5D4(
.data_in(MC_L1L2_L5D4_FM_L1L2_L5D4),
.enable(MC_L1L2_L5D4_FM_L1L2_L5D4_wr_en),
.number_out(FM_L1L2_L5D4_FT_L1L2_number),
.read_add(FM_L1L2_L5D4_FT_L1L2_read_add),
.data_out(FM_L1L2_L5D4_FT_L1L2),
.read_en(FM_L1L2_L5D4_FT_L1L2_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L6D3_FM_L1L2_L6D3;
wire MC_L1L2_L6D3_FM_L1L2_L6D3_wr_en;
wire [5:0] FM_L1L2_L6D3_FT_L1L2_number;
wire [9:0] FM_L1L2_L6D3_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L6D3_FT_L1L2;
wire FM_L1L2_L6D3_FT_L1L2_read_en;
FullMatch  FM_L1L2_L6D3(
.data_in(MC_L1L2_L6D3_FM_L1L2_L6D3),
.enable(MC_L1L2_L6D3_FM_L1L2_L6D3_wr_en),
.number_out(FM_L1L2_L6D3_FT_L1L2_number),
.read_add(FM_L1L2_L6D3_FT_L1L2_read_add),
.data_out(FM_L1L2_L6D3_FT_L1L2),
.read_en(FM_L1L2_L6D3_FT_L1L2_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L1L2_L6D4_FM_L1L2_L6D4;
wire MC_L1L2_L6D4_FM_L1L2_L6D4_wr_en;
wire [5:0] FM_L1L2_L6D4_FT_L1L2_number;
wire [9:0] FM_L1L2_L6D4_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L6D4_FT_L1L2;
wire FM_L1L2_L6D4_FT_L1L2_read_en;
FullMatch  FM_L1L2_L6D4(
.data_in(MC_L1L2_L6D4_FM_L1L2_L6D4),
.enable(MC_L1L2_L6D4_FM_L1L2_L6D4_wr_en),
.number_out(FM_L1L2_L6D4_FT_L1L2_number),
.read_add(FM_L1L2_L6D4_FT_L1L2_read_add),
.data_out(FM_L1L2_L6D4_FT_L1L2),
.read_en(FM_L1L2_L6D4_FT_L1L2_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L1D3L2D3_TPAR_L1D3L2D3;
wire TC_L1D3L2D3_TPAR_L1D3L2D3_wr_en;
wire [10:0] TPAR_L1D3L2D3_FT_L1L2_read_add;
wire [55:0] TPAR_L1D3L2D3_FT_L1L2;
TrackletParameters  TPAR_L1D3L2D3(
.data_in(TC_L1D3L2D3_TPAR_L1D3L2D3),
.enable(TC_L1D3L2D3_TPAR_L1D3L2D3_wr_en),
.read_add(TPAR_L1D3L2D3_FT_L1L2_read_add),
.data_out(TPAR_L1D3L2D3_FT_L1L2),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L1D3L2D4_TPAR_L1D3L2D4;
wire TC_L1D3L2D4_TPAR_L1D3L2D4_wr_en;
wire [10:0] TPAR_L1D3L2D4_FT_L1L2_read_add;
wire [55:0] TPAR_L1D3L2D4_FT_L1L2;
TrackletParameters  TPAR_L1D3L2D4(
.data_in(TC_L1D3L2D4_TPAR_L1D3L2D4),
.enable(TC_L1D3L2D4_TPAR_L1D3L2D4_wr_en),
.read_add(TPAR_L1D3L2D4_FT_L1L2_read_add),
.data_out(TPAR_L1D3L2D4_FT_L1L2),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L1D4L2D4_TPAR_L1D4L2D4;
wire TC_L1D4L2D4_TPAR_L1D4L2D4_wr_en;
wire [10:0] TPAR_L1D4L2D4_FT_L1L2_read_add;
wire [55:0] TPAR_L1D4L2D4_FT_L1L2;
TrackletParameters  TPAR_L1D4L2D4(
.data_in(TC_L1D4L2D4_TPAR_L1D4L2D4),
.enable(TC_L1D4L2D4_TPAR_L1D4L2D4_wr_en),
.read_add(TPAR_L1D4L2D4_FT_L1L2_read_add),
.data_out(TPAR_L1D4L2D4_FT_L1L2),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L1L2_Plus_FM_L1L2_L3_FromPlus;
wire MT_L1L2_Plus_FM_L1L2_L3_FromPlus_wr_en;
wire [5:0] FM_L1L2_L3_FromPlus_FT_L1L2_number;
wire [9:0] FM_L1L2_L3_FromPlus_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L3_FromPlus_FT_L1L2;
wire FM_L1L2_L3_FromPlus_FT_L1L2_read_en;
FullMatch #(128) FM_L1L2_L3_FromPlus(
.data_in(MT_L1L2_Plus_FM_L1L2_L3_FromPlus),
.enable(MT_L1L2_Plus_FM_L1L2_L3_FromPlus_wr_en),
.number_out(FM_L1L2_L3_FromPlus_FT_L1L2_number),
.read_add(FM_L1L2_L3_FromPlus_FT_L1L2_read_add),
.data_out(FM_L1L2_L3_FromPlus_FT_L1L2),
.read_en(FM_L1L2_L3_FromPlus_FT_L1L2_read_en),
.start(start10_0),
.done(done9_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L1L2_Plus_FM_L1L2_L4_FromPlus;
wire MT_L1L2_Plus_FM_L1L2_L4_FromPlus_wr_en;
wire [5:0] FM_L1L2_L4_FromPlus_FT_L1L2_number;
wire [9:0] FM_L1L2_L4_FromPlus_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L4_FromPlus_FT_L1L2;
wire FM_L1L2_L4_FromPlus_FT_L1L2_read_en;
FullMatch #(128) FM_L1L2_L4_FromPlus(
.data_in(MT_L1L2_Plus_FM_L1L2_L4_FromPlus),
.enable(MT_L1L2_Plus_FM_L1L2_L4_FromPlus_wr_en),
.number_out(FM_L1L2_L4_FromPlus_FT_L1L2_number),
.read_add(FM_L1L2_L4_FromPlus_FT_L1L2_read_add),
.data_out(FM_L1L2_L4_FromPlus_FT_L1L2),
.read_en(FM_L1L2_L4_FromPlus_FT_L1L2_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L1L2_Plus_FM_L1L2_L5_FromPlus;
wire MT_L1L2_Plus_FM_L1L2_L5_FromPlus_wr_en;
wire [5:0] FM_L1L2_L5_FromPlus_FT_L1L2_number;
wire [9:0] FM_L1L2_L5_FromPlus_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L5_FromPlus_FT_L1L2;
wire FM_L1L2_L5_FromPlus_FT_L1L2_read_en;
FullMatch #(128) FM_L1L2_L5_FromPlus(
.data_in(MT_L1L2_Plus_FM_L1L2_L5_FromPlus),
.enable(MT_L1L2_Plus_FM_L1L2_L5_FromPlus_wr_en),
.number_out(FM_L1L2_L5_FromPlus_FT_L1L2_number),
.read_add(FM_L1L2_L5_FromPlus_FT_L1L2_read_add),
.data_out(FM_L1L2_L5_FromPlus_FT_L1L2),
.read_en(FM_L1L2_L5_FromPlus_FT_L1L2_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L1L2_Plus_FM_L1L2_L6_FromPlus;
wire MT_L1L2_Plus_FM_L1L2_L6_FromPlus_wr_en;
wire [5:0] FM_L1L2_L6_FromPlus_FT_L1L2_number;
wire [9:0] FM_L1L2_L6_FromPlus_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L6_FromPlus_FT_L1L2;
wire FM_L1L2_L6_FromPlus_FT_L1L2_read_en;
FullMatch #(128) FM_L1L2_L6_FromPlus(
.data_in(MT_L1L2_Plus_FM_L1L2_L6_FromPlus),
.enable(MT_L1L2_Plus_FM_L1L2_L6_FromPlus_wr_en),
.number_out(FM_L1L2_L6_FromPlus_FT_L1L2_number),
.read_add(FM_L1L2_L6_FromPlus_FT_L1L2_read_add),
.data_out(FM_L1L2_L6_FromPlus_FT_L1L2),
.read_en(FM_L1L2_L6_FromPlus_FT_L1L2_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L1L2_Minus_FM_L1L2_L3_FromMinus;
wire MT_L1L2_Minus_FM_L1L2_L3_FromMinus_wr_en;
wire [5:0] FM_L1L2_L3_FromMinus_FT_L1L2_number;
wire [9:0] FM_L1L2_L3_FromMinus_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L3_FromMinus_FT_L1L2;
wire FM_L1L2_L3_FromMinus_FT_L1L2_read_en;
FullMatch #(128) FM_L1L2_L3_FromMinus(
.data_in(MT_L1L2_Minus_FM_L1L2_L3_FromMinus),
.enable(MT_L1L2_Minus_FM_L1L2_L3_FromMinus_wr_en),
.number_out(FM_L1L2_L3_FromMinus_FT_L1L2_number),
.read_add(FM_L1L2_L3_FromMinus_FT_L1L2_read_add),
.data_out(FM_L1L2_L3_FromMinus_FT_L1L2),
.read_en(FM_L1L2_L3_FromMinus_FT_L1L2_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L1L2_Minus_FM_L1L2_L4_FromMinus;
wire MT_L1L2_Minus_FM_L1L2_L4_FromMinus_wr_en;
wire [5:0] FM_L1L2_L4_FromMinus_FT_L1L2_number;
wire [9:0] FM_L1L2_L4_FromMinus_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L4_FromMinus_FT_L1L2;
wire FM_L1L2_L4_FromMinus_FT_L1L2_read_en;
FullMatch #(128) FM_L1L2_L4_FromMinus(
.data_in(MT_L1L2_Minus_FM_L1L2_L4_FromMinus),
.enable(MT_L1L2_Minus_FM_L1L2_L4_FromMinus_wr_en),
.number_out(FM_L1L2_L4_FromMinus_FT_L1L2_number),
.read_add(FM_L1L2_L4_FromMinus_FT_L1L2_read_add),
.data_out(FM_L1L2_L4_FromMinus_FT_L1L2),
.read_en(FM_L1L2_L4_FromMinus_FT_L1L2_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L1L2_Minus_FM_L1L2_L5_FromMinus;
wire MT_L1L2_Minus_FM_L1L2_L5_FromMinus_wr_en;
wire [5:0] FM_L1L2_L5_FromMinus_FT_L1L2_number;
wire [9:0] FM_L1L2_L5_FromMinus_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L5_FromMinus_FT_L1L2;
wire FM_L1L2_L5_FromMinus_FT_L1L2_read_en;
FullMatch #(128) FM_L1L2_L5_FromMinus(
.data_in(MT_L1L2_Minus_FM_L1L2_L5_FromMinus),
.enable(MT_L1L2_Minus_FM_L1L2_L5_FromMinus_wr_en),
.number_out(FM_L1L2_L5_FromMinus_FT_L1L2_number),
.read_add(FM_L1L2_L5_FromMinus_FT_L1L2_read_add),
.data_out(FM_L1L2_L5_FromMinus_FT_L1L2),
.read_en(FM_L1L2_L5_FromMinus_FT_L1L2_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L1L2_Minus_FM_L1L2_L6_FromMinus;
wire MT_L1L2_Minus_FM_L1L2_L6_FromMinus_wr_en;
wire [5:0] FM_L1L2_L6_FromMinus_FT_L1L2_number;
wire [9:0] FM_L1L2_L6_FromMinus_FT_L1L2_read_add;
wire [35:0] FM_L1L2_L6_FromMinus_FT_L1L2;
wire FM_L1L2_L6_FromMinus_FT_L1L2_read_en;
FullMatch #(128) FM_L1L2_L6_FromMinus(
.data_in(MT_L1L2_Minus_FM_L1L2_L6_FromMinus),
.enable(MT_L1L2_Minus_FM_L1L2_L6_FromMinus_wr_en),
.number_out(FM_L1L2_L6_FromMinus_FT_L1L2_number),
.read_add(FM_L1L2_L6_FromMinus_FT_L1L2_read_add),
.data_out(FM_L1L2_L6_FromMinus_FT_L1L2),
.read_en(FM_L1L2_L6_FromMinus_FT_L1L2_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L1D3_FM_L3L4_L1D3;
wire MC_L3L4_L1D3_FM_L3L4_L1D3_wr_en;
wire [5:0] FM_L3L4_L1D3_FT_L3L4_number;
wire [9:0] FM_L3L4_L1D3_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L1D3_FT_L3L4;
wire FM_L3L4_L1D3_FT_L3L4_read_en;
FullMatch  FM_L3L4_L1D3(
.data_in(MC_L3L4_L1D3_FM_L3L4_L1D3),
.enable(MC_L3L4_L1D3_FM_L3L4_L1D3_wr_en),
.number_out(FM_L3L4_L1D3_FT_L3L4_number),
.read_add(FM_L3L4_L1D3_FT_L3L4_read_add),
.data_out(FM_L3L4_L1D3_FT_L3L4),
.read_en(FM_L3L4_L1D3_FT_L3L4_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L1D4_FM_L3L4_L1D4;
wire MC_L3L4_L1D4_FM_L3L4_L1D4_wr_en;
wire [5:0] FM_L3L4_L1D4_FT_L3L4_number;
wire [9:0] FM_L3L4_L1D4_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L1D4_FT_L3L4;
wire FM_L3L4_L1D4_FT_L3L4_read_en;
FullMatch  FM_L3L4_L1D4(
.data_in(MC_L3L4_L1D4_FM_L3L4_L1D4),
.enable(MC_L3L4_L1D4_FM_L3L4_L1D4_wr_en),
.number_out(FM_L3L4_L1D4_FT_L3L4_number),
.read_add(FM_L3L4_L1D4_FT_L3L4_read_add),
.data_out(FM_L3L4_L1D4_FT_L3L4),
.read_en(FM_L3L4_L1D4_FT_L3L4_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L2D3_FM_L3L4_L2D3;
wire MC_L3L4_L2D3_FM_L3L4_L2D3_wr_en;
wire [5:0] FM_L3L4_L2D3_FT_L3L4_number;
wire [9:0] FM_L3L4_L2D3_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L2D3_FT_L3L4;
wire FM_L3L4_L2D3_FT_L3L4_read_en;
FullMatch  FM_L3L4_L2D3(
.data_in(MC_L3L4_L2D3_FM_L3L4_L2D3),
.enable(MC_L3L4_L2D3_FM_L3L4_L2D3_wr_en),
.number_out(FM_L3L4_L2D3_FT_L3L4_number),
.read_add(FM_L3L4_L2D3_FT_L3L4_read_add),
.data_out(FM_L3L4_L2D3_FT_L3L4),
.read_en(FM_L3L4_L2D3_FT_L3L4_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L2D4_FM_L3L4_L2D4;
wire MC_L3L4_L2D4_FM_L3L4_L2D4_wr_en;
wire [5:0] FM_L3L4_L2D4_FT_L3L4_number;
wire [9:0] FM_L3L4_L2D4_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L2D4_FT_L3L4;
wire FM_L3L4_L2D4_FT_L3L4_read_en;
FullMatch  FM_L3L4_L2D4(
.data_in(MC_L3L4_L2D4_FM_L3L4_L2D4),
.enable(MC_L3L4_L2D4_FM_L3L4_L2D4_wr_en),
.number_out(FM_L3L4_L2D4_FT_L3L4_number),
.read_add(FM_L3L4_L2D4_FT_L3L4_read_add),
.data_out(FM_L3L4_L2D4_FT_L3L4),
.read_en(FM_L3L4_L2D4_FT_L3L4_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L5D3_FM_L3L4_L5D3;
wire MC_L3L4_L5D3_FM_L3L4_L5D3_wr_en;
wire [5:0] FM_L3L4_L5D3_FT_L3L4_number;
wire [9:0] FM_L3L4_L5D3_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L5D3_FT_L3L4;
wire FM_L3L4_L5D3_FT_L3L4_read_en;
FullMatch  FM_L3L4_L5D3(
.data_in(MC_L3L4_L5D3_FM_L3L4_L5D3),
.enable(MC_L3L4_L5D3_FM_L3L4_L5D3_wr_en),
.number_out(FM_L3L4_L5D3_FT_L3L4_number),
.read_add(FM_L3L4_L5D3_FT_L3L4_read_add),
.data_out(FM_L3L4_L5D3_FT_L3L4),
.read_en(FM_L3L4_L5D3_FT_L3L4_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L5D4_FM_L3L4_L5D4;
wire MC_L3L4_L5D4_FM_L3L4_L5D4_wr_en;
wire [5:0] FM_L3L4_L5D4_FT_L3L4_number;
wire [9:0] FM_L3L4_L5D4_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L5D4_FT_L3L4;
wire FM_L3L4_L5D4_FT_L3L4_read_en;
FullMatch  FM_L3L4_L5D4(
.data_in(MC_L3L4_L5D4_FM_L3L4_L5D4),
.enable(MC_L3L4_L5D4_FM_L3L4_L5D4_wr_en),
.number_out(FM_L3L4_L5D4_FT_L3L4_number),
.read_add(FM_L3L4_L5D4_FT_L3L4_read_add),
.data_out(FM_L3L4_L5D4_FT_L3L4),
.read_en(FM_L3L4_L5D4_FT_L3L4_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L6D3_FM_L3L4_L6D3;
wire MC_L3L4_L6D3_FM_L3L4_L6D3_wr_en;
wire [5:0] FM_L3L4_L6D3_FT_L3L4_number;
wire [9:0] FM_L3L4_L6D3_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L6D3_FT_L3L4;
wire FM_L3L4_L6D3_FT_L3L4_read_en;
FullMatch  FM_L3L4_L6D3(
.data_in(MC_L3L4_L6D3_FM_L3L4_L6D3),
.enable(MC_L3L4_L6D3_FM_L3L4_L6D3_wr_en),
.number_out(FM_L3L4_L6D3_FT_L3L4_number),
.read_add(FM_L3L4_L6D3_FT_L3L4_read_add),
.data_out(FM_L3L4_L6D3_FT_L3L4),
.read_en(FM_L3L4_L6D3_FT_L3L4_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L3L4_L6D4_FM_L3L4_L6D4;
wire MC_L3L4_L6D4_FM_L3L4_L6D4_wr_en;
wire [5:0] FM_L3L4_L6D4_FT_L3L4_number;
wire [9:0] FM_L3L4_L6D4_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L6D4_FT_L3L4;
wire FM_L3L4_L6D4_FT_L3L4_read_en;
FullMatch  FM_L3L4_L6D4(
.data_in(MC_L3L4_L6D4_FM_L3L4_L6D4),
.enable(MC_L3L4_L6D4_FM_L3L4_L6D4_wr_en),
.number_out(FM_L3L4_L6D4_FT_L3L4_number),
.read_add(FM_L3L4_L6D4_FT_L3L4_read_add),
.data_out(FM_L3L4_L6D4_FT_L3L4),
.read_en(FM_L3L4_L6D4_FT_L3L4_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L3L4_Minus_FM_L3L4_L1_FromMinus;
wire MT_L3L4_Minus_FM_L3L4_L1_FromMinus_wr_en;
wire [5:0] FM_L3L4_L1_FromMinus_FT_L3L4_number;
wire [9:0] FM_L3L4_L1_FromMinus_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L1_FromMinus_FT_L3L4;
wire FM_L3L4_L1_FromMinus_FT_L3L4_read_en;
FullMatch #(128) FM_L3L4_L1_FromMinus(
.data_in(MT_L3L4_Minus_FM_L3L4_L1_FromMinus),
.enable(MT_L3L4_Minus_FM_L3L4_L1_FromMinus_wr_en),
.number_out(FM_L3L4_L1_FromMinus_FT_L3L4_number),
.read_add(FM_L3L4_L1_FromMinus_FT_L3L4_read_add),
.data_out(FM_L3L4_L1_FromMinus_FT_L3L4),
.read_en(FM_L3L4_L1_FromMinus_FT_L3L4_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L3L4_Minus_FM_L3L4_L2_FromMinus;
wire MT_L3L4_Minus_FM_L3L4_L2_FromMinus_wr_en;
wire [5:0] FM_L3L4_L2_FromMinus_FT_L3L4_number;
wire [9:0] FM_L3L4_L2_FromMinus_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L2_FromMinus_FT_L3L4;
wire FM_L3L4_L2_FromMinus_FT_L3L4_read_en;
FullMatch #(128) FM_L3L4_L2_FromMinus(
.data_in(MT_L3L4_Minus_FM_L3L4_L2_FromMinus),
.enable(MT_L3L4_Minus_FM_L3L4_L2_FromMinus_wr_en),
.number_out(FM_L3L4_L2_FromMinus_FT_L3L4_number),
.read_add(FM_L3L4_L2_FromMinus_FT_L3L4_read_add),
.data_out(FM_L3L4_L2_FromMinus_FT_L3L4),
.read_en(FM_L3L4_L2_FromMinus_FT_L3L4_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L3L4_Minus_FM_L3L4_L5_FromMinus;
wire MT_L3L4_Minus_FM_L3L4_L5_FromMinus_wr_en;
wire [5:0] FM_L3L4_L5_FromMinus_FT_L3L4_number;
wire [9:0] FM_L3L4_L5_FromMinus_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L5_FromMinus_FT_L3L4;
wire FM_L3L4_L5_FromMinus_FT_L3L4_read_en;
FullMatch #(128) FM_L3L4_L5_FromMinus(
.data_in(MT_L3L4_Minus_FM_L3L4_L5_FromMinus),
.enable(MT_L3L4_Minus_FM_L3L4_L5_FromMinus_wr_en),
.number_out(FM_L3L4_L5_FromMinus_FT_L3L4_number),
.read_add(FM_L3L4_L5_FromMinus_FT_L3L4_read_add),
.data_out(FM_L3L4_L5_FromMinus_FT_L3L4),
.read_en(FM_L3L4_L5_FromMinus_FT_L3L4_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L3L4_Minus_FM_L3L4_L6_FromMinus;
wire MT_L3L4_Minus_FM_L3L4_L6_FromMinus_wr_en;
wire [5:0] FM_L3L4_L6_FromMinus_FT_L3L4_number;
wire [9:0] FM_L3L4_L6_FromMinus_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L6_FromMinus_FT_L3L4;
wire FM_L3L4_L6_FromMinus_FT_L3L4_read_en;
FullMatch #(128) FM_L3L4_L6_FromMinus(
.data_in(MT_L3L4_Minus_FM_L3L4_L6_FromMinus),
.enable(MT_L3L4_Minus_FM_L3L4_L6_FromMinus_wr_en),
.number_out(FM_L3L4_L6_FromMinus_FT_L3L4_number),
.read_add(FM_L3L4_L6_FromMinus_FT_L3L4_read_add),
.data_out(FM_L3L4_L6_FromMinus_FT_L3L4),
.read_en(FM_L3L4_L6_FromMinus_FT_L3L4_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L3L4_Plus_FM_L3L4_L1_FromPlus;
wire MT_L3L4_Plus_FM_L3L4_L1_FromPlus_wr_en;
wire [5:0] FM_L3L4_L1_FromPlus_FT_L3L4_number;
wire [9:0] FM_L3L4_L1_FromPlus_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L1_FromPlus_FT_L3L4;
wire FM_L3L4_L1_FromPlus_FT_L3L4_read_en;
FullMatch #(128) FM_L3L4_L1_FromPlus(
.data_in(MT_L3L4_Plus_FM_L3L4_L1_FromPlus),
.enable(MT_L3L4_Plus_FM_L3L4_L1_FromPlus_wr_en),
.number_out(FM_L3L4_L1_FromPlus_FT_L3L4_number),
.read_add(FM_L3L4_L1_FromPlus_FT_L3L4_read_add),
.data_out(FM_L3L4_L1_FromPlus_FT_L3L4),
.read_en(FM_L3L4_L1_FromPlus_FT_L3L4_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L3L4_Plus_FM_L3L4_L2_FromPlus;
wire MT_L3L4_Plus_FM_L3L4_L2_FromPlus_wr_en;
wire [5:0] FM_L3L4_L2_FromPlus_FT_L3L4_number;
wire [9:0] FM_L3L4_L2_FromPlus_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L2_FromPlus_FT_L3L4;
wire FM_L3L4_L2_FromPlus_FT_L3L4_read_en;
FullMatch #(128) FM_L3L4_L2_FromPlus(
.data_in(MT_L3L4_Plus_FM_L3L4_L2_FromPlus),
.enable(MT_L3L4_Plus_FM_L3L4_L2_FromPlus_wr_en),
.number_out(FM_L3L4_L2_FromPlus_FT_L3L4_number),
.read_add(FM_L3L4_L2_FromPlus_FT_L3L4_read_add),
.data_out(FM_L3L4_L2_FromPlus_FT_L3L4),
.read_en(FM_L3L4_L2_FromPlus_FT_L3L4_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L3L4_Plus_FM_L3L4_L5_FromPlus;
wire MT_L3L4_Plus_FM_L3L4_L5_FromPlus_wr_en;
wire [5:0] FM_L3L4_L5_FromPlus_FT_L3L4_number;
wire [9:0] FM_L3L4_L5_FromPlus_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L5_FromPlus_FT_L3L4;
wire FM_L3L4_L5_FromPlus_FT_L3L4_read_en;
FullMatch #(128) FM_L3L4_L5_FromPlus(
.data_in(MT_L3L4_Plus_FM_L3L4_L5_FromPlus),
.enable(MT_L3L4_Plus_FM_L3L4_L5_FromPlus_wr_en),
.number_out(FM_L3L4_L5_FromPlus_FT_L3L4_number),
.read_add(FM_L3L4_L5_FromPlus_FT_L3L4_read_add),
.data_out(FM_L3L4_L5_FromPlus_FT_L3L4),
.read_en(FM_L3L4_L5_FromPlus_FT_L3L4_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L3L4_Plus_FM_L3L4_L6_FromPlus;
wire MT_L3L4_Plus_FM_L3L4_L6_FromPlus_wr_en;
wire [5:0] FM_L3L4_L6_FromPlus_FT_L3L4_number;
wire [9:0] FM_L3L4_L6_FromPlus_FT_L3L4_read_add;
wire [35:0] FM_L3L4_L6_FromPlus_FT_L3L4;
wire FM_L3L4_L6_FromPlus_FT_L3L4_read_en;
FullMatch #(128) FM_L3L4_L6_FromPlus(
.data_in(MT_L3L4_Plus_FM_L3L4_L6_FromPlus),
.enable(MT_L3L4_Plus_FM_L3L4_L6_FromPlus_wr_en),
.number_out(FM_L3L4_L6_FromPlus_FT_L3L4_number),
.read_add(FM_L3L4_L6_FromPlus_FT_L3L4_read_add),
.data_out(FM_L3L4_L6_FromPlus_FT_L3L4),
.read_en(FM_L3L4_L6_FromPlus_FT_L3L4_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L3D3L4D3_TPAR_L3D3L4D3;
wire TC_L3D3L4D3_TPAR_L3D3L4D3_wr_en;
wire [10:0] TPAR_L3D3L4D3_FT_L3L4_read_add;
wire [55:0] TPAR_L3D3L4D3_FT_L3L4;
TrackletParameters  TPAR_L3D3L4D3(
.data_in(TC_L3D3L4D3_TPAR_L3D3L4D3),
.enable(TC_L3D3L4D3_TPAR_L3D3L4D3_wr_en),
.read_add(TPAR_L3D3L4D3_FT_L3L4_read_add),
.data_out(TPAR_L3D3L4D3_FT_L3L4),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L3D3L4D4_TPAR_L3D3L4D4;
wire TC_L3D3L4D4_TPAR_L3D3L4D4_wr_en;
wire [10:0] TPAR_L3D3L4D4_FT_L3L4_read_add;
wire [55:0] TPAR_L3D3L4D4_FT_L3L4;
TrackletParameters  TPAR_L3D3L4D4(
.data_in(TC_L3D3L4D4_TPAR_L3D3L4D4),
.enable(TC_L3D3L4D4_TPAR_L3D3L4D4_wr_en),
.read_add(TPAR_L3D3L4D4_FT_L3L4_read_add),
.data_out(TPAR_L3D3L4D4_FT_L3L4),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L3D4L4D4_TPAR_L3D4L4D4;
wire TC_L3D4L4D4_TPAR_L3D4L4D4_wr_en;
wire [10:0] TPAR_L3D4L4D4_FT_L3L4_read_add;
wire [55:0] TPAR_L3D4L4D4_FT_L3L4;
TrackletParameters  TPAR_L3D4L4D4(
.data_in(TC_L3D4L4D4_TPAR_L3D4L4D4),
.enable(TC_L3D4L4D4_TPAR_L3D4L4D4_wr_en),
.read_add(TPAR_L3D4L4D4_FT_L3L4_read_add),
.data_out(TPAR_L3D4L4D4_FT_L3L4),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L1D3_FM_L5L6_L1D3;
wire MC_L5L6_L1D3_FM_L5L6_L1D3_wr_en;
wire [5:0] FM_L5L6_L1D3_FT_L5L6_number;
wire [9:0] FM_L5L6_L1D3_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L1D3_FT_L5L6;
wire FM_L5L6_L1D3_FT_L5L6_read_en;
FullMatch  FM_L5L6_L1D3(
.data_in(MC_L5L6_L1D3_FM_L5L6_L1D3),
.enable(MC_L5L6_L1D3_FM_L5L6_L1D3_wr_en),
.number_out(FM_L5L6_L1D3_FT_L5L6_number),
.read_add(FM_L5L6_L1D3_FT_L5L6_read_add),
.data_out(FM_L5L6_L1D3_FT_L5L6),
.read_en(FM_L5L6_L1D3_FT_L5L6_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L1D4_FM_L5L6_L1D4;
wire MC_L5L6_L1D4_FM_L5L6_L1D4_wr_en;
wire [5:0] FM_L5L6_L1D4_FT_L5L6_number;
wire [9:0] FM_L5L6_L1D4_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L1D4_FT_L5L6;
wire FM_L5L6_L1D4_FT_L5L6_read_en;
FullMatch  FM_L5L6_L1D4(
.data_in(MC_L5L6_L1D4_FM_L5L6_L1D4),
.enable(MC_L5L6_L1D4_FM_L5L6_L1D4_wr_en),
.number_out(FM_L5L6_L1D4_FT_L5L6_number),
.read_add(FM_L5L6_L1D4_FT_L5L6_read_add),
.data_out(FM_L5L6_L1D4_FT_L5L6),
.read_en(FM_L5L6_L1D4_FT_L5L6_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L2D3_FM_L5L6_L2D3;
wire MC_L5L6_L2D3_FM_L5L6_L2D3_wr_en;
wire [5:0] FM_L5L6_L2D3_FT_L5L6_number;
wire [9:0] FM_L5L6_L2D3_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L2D3_FT_L5L6;
wire FM_L5L6_L2D3_FT_L5L6_read_en;
FullMatch  FM_L5L6_L2D3(
.data_in(MC_L5L6_L2D3_FM_L5L6_L2D3),
.enable(MC_L5L6_L2D3_FM_L5L6_L2D3_wr_en),
.number_out(FM_L5L6_L2D3_FT_L5L6_number),
.read_add(FM_L5L6_L2D3_FT_L5L6_read_add),
.data_out(FM_L5L6_L2D3_FT_L5L6),
.read_en(FM_L5L6_L2D3_FT_L5L6_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L2D4_FM_L5L6_L2D4;
wire MC_L5L6_L2D4_FM_L5L6_L2D4_wr_en;
wire [5:0] FM_L5L6_L2D4_FT_L5L6_number;
wire [9:0] FM_L5L6_L2D4_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L2D4_FT_L5L6;
wire FM_L5L6_L2D4_FT_L5L6_read_en;
FullMatch  FM_L5L6_L2D4(
.data_in(MC_L5L6_L2D4_FM_L5L6_L2D4),
.enable(MC_L5L6_L2D4_FM_L5L6_L2D4_wr_en),
.number_out(FM_L5L6_L2D4_FT_L5L6_number),
.read_add(FM_L5L6_L2D4_FT_L5L6_read_add),
.data_out(FM_L5L6_L2D4_FT_L5L6),
.read_en(FM_L5L6_L2D4_FT_L5L6_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L3D3_FM_L5L6_L3D3;
wire MC_L5L6_L3D3_FM_L5L6_L3D3_wr_en;
wire [5:0] FM_L5L6_L3D3_FT_L5L6_number;
wire [9:0] FM_L5L6_L3D3_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L3D3_FT_L5L6;
wire FM_L5L6_L3D3_FT_L5L6_read_en;
FullMatch  FM_L5L6_L3D3(
.data_in(MC_L5L6_L3D3_FM_L5L6_L3D3),
.enable(MC_L5L6_L3D3_FM_L5L6_L3D3_wr_en),
.number_out(FM_L5L6_L3D3_FT_L5L6_number),
.read_add(FM_L5L6_L3D3_FT_L5L6_read_add),
.data_out(FM_L5L6_L3D3_FT_L5L6),
.read_en(FM_L5L6_L3D3_FT_L5L6_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L3D4_FM_L5L6_L3D4;
wire MC_L5L6_L3D4_FM_L5L6_L3D4_wr_en;
wire [5:0] FM_L5L6_L3D4_FT_L5L6_number;
wire [9:0] FM_L5L6_L3D4_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L3D4_FT_L5L6;
wire FM_L5L6_L3D4_FT_L5L6_read_en;
FullMatch  FM_L5L6_L3D4(
.data_in(MC_L5L6_L3D4_FM_L5L6_L3D4),
.enable(MC_L5L6_L3D4_FM_L5L6_L3D4_wr_en),
.number_out(FM_L5L6_L3D4_FT_L5L6_number),
.read_add(FM_L5L6_L3D4_FT_L5L6_read_add),
.data_out(FM_L5L6_L3D4_FT_L5L6),
.read_en(FM_L5L6_L3D4_FT_L5L6_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L4D3_FM_L5L6_L4D3;
wire MC_L5L6_L4D3_FM_L5L6_L4D3_wr_en;
wire [5:0] FM_L5L6_L4D3_FT_L5L6_number;
wire [9:0] FM_L5L6_L4D3_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L4D3_FT_L5L6;
wire FM_L5L6_L4D3_FT_L5L6_read_en;
FullMatch  FM_L5L6_L4D3(
.data_in(MC_L5L6_L4D3_FM_L5L6_L4D3),
.enable(MC_L5L6_L4D3_FM_L5L6_L4D3_wr_en),
.number_out(FM_L5L6_L4D3_FT_L5L6_number),
.read_add(FM_L5L6_L4D3_FT_L5L6_read_add),
.data_out(FM_L5L6_L4D3_FT_L5L6),
.read_en(FM_L5L6_L4D3_FT_L5L6_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MC_L5L6_L4D4_FM_L5L6_L4D4;
wire MC_L5L6_L4D4_FM_L5L6_L4D4_wr_en;
wire [5:0] FM_L5L6_L4D4_FT_L5L6_number;
wire [9:0] FM_L5L6_L4D4_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L4D4_FT_L5L6;
wire FM_L5L6_L4D4_FT_L5L6_read_en;
FullMatch  FM_L5L6_L4D4(
.data_in(MC_L5L6_L4D4_FM_L5L6_L4D4),
.enable(MC_L5L6_L4D4_FM_L5L6_L4D4_wr_en),
.number_out(FM_L5L6_L4D4_FT_L5L6_number),
.read_add(FM_L5L6_L4D4_FT_L5L6_read_add),
.data_out(FM_L5L6_L4D4_FT_L5L6),
.read_en(FM_L5L6_L4D4_FT_L5L6_read_en),
.start(start9_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L5D3L6D3_TPAR_L5D3L6D3;
wire TC_L5D3L6D3_TPAR_L5D3L6D3_wr_en;
wire [10:0] TPAR_L5D3L6D3_FT_L5L6_read_add;
wire [55:0] TPAR_L5D3L6D3_FT_L5L6;
TrackletParameters  TPAR_L5D3L6D3(
.data_in(TC_L5D3L6D3_TPAR_L5D3L6D3),
.enable(TC_L5D3L6D3_TPAR_L5D3L6D3_wr_en),
.read_add(TPAR_L5D3L6D3_FT_L5L6_read_add),
.data_out(TPAR_L5D3L6D3_FT_L5L6),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L5D3L6D4_TPAR_L5D3L6D4;
wire TC_L5D3L6D4_TPAR_L5D3L6D4_wr_en;
wire [10:0] TPAR_L5D3L6D4_FT_L5L6_read_add;
wire [55:0] TPAR_L5D3L6D4_FT_L5L6;
TrackletParameters  TPAR_L5D3L6D4(
.data_in(TC_L5D3L6D4_TPAR_L5D3L6D4),
.enable(TC_L5D3L6D4_TPAR_L5D3L6D4_wr_en),
.read_add(TPAR_L5D3L6D4_FT_L5L6_read_add),
.data_out(TPAR_L5D3L6D4_FT_L5L6),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [55:0] TC_L5D4L6D4_TPAR_L5D4L6D4;
wire TC_L5D4L6D4_TPAR_L5D4L6D4_wr_en;
wire [10:0] TPAR_L5D4L6D4_FT_L5L6_read_add;
wire [55:0] TPAR_L5D4L6D4_FT_L5L6;
TrackletParameters  TPAR_L5D4L6D4(
.data_in(TC_L5D4L6D4_TPAR_L5D4L6D4),
.enable(TC_L5D4L6D4_TPAR_L5D4L6D4_wr_en),
.read_add(TPAR_L5D4L6D4_FT_L5L6_read_add),
.data_out(TPAR_L5D4L6D4_FT_L5L6),
.start(start5_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L5L6_Plus_FM_L5L6_L1_FromPlus;
wire MT_L5L6_Plus_FM_L5L6_L1_FromPlus_wr_en;
wire [5:0] FM_L5L6_L1_FromPlus_FT_L5L6_number;
wire [9:0] FM_L5L6_L1_FromPlus_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L1_FromPlus_FT_L5L6;
wire FM_L5L6_L1_FromPlus_FT_L5L6_read_en;
FullMatch #(128) FM_L5L6_L1_FromPlus(
.data_in(MT_L5L6_Plus_FM_L5L6_L1_FromPlus),
.enable(MT_L5L6_Plus_FM_L5L6_L1_FromPlus_wr_en),
.number_out(FM_L5L6_L1_FromPlus_FT_L5L6_number),
.read_add(FM_L5L6_L1_FromPlus_FT_L5L6_read_add),
.data_out(FM_L5L6_L1_FromPlus_FT_L5L6),
.read_en(FM_L5L6_L1_FromPlus_FT_L5L6_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L5L6_Plus_FM_L5L6_L2_FromPlus;
wire MT_L5L6_Plus_FM_L5L6_L2_FromPlus_wr_en;
wire [5:0] FM_L5L6_L2_FromPlus_FT_L5L6_number;
wire [9:0] FM_L5L6_L2_FromPlus_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L2_FromPlus_FT_L5L6;
wire FM_L5L6_L2_FromPlus_FT_L5L6_read_en;
FullMatch #(128) FM_L5L6_L2_FromPlus(
.data_in(MT_L5L6_Plus_FM_L5L6_L2_FromPlus),
.enable(MT_L5L6_Plus_FM_L5L6_L2_FromPlus_wr_en),
.number_out(FM_L5L6_L2_FromPlus_FT_L5L6_number),
.read_add(FM_L5L6_L2_FromPlus_FT_L5L6_read_add),
.data_out(FM_L5L6_L2_FromPlus_FT_L5L6),
.read_en(FM_L5L6_L2_FromPlus_FT_L5L6_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L5L6_Plus_FM_L5L6_L3_FromPlus;
wire MT_L5L6_Plus_FM_L5L6_L3_FromPlus_wr_en;
wire [5:0] FM_L5L6_L3_FromPlus_FT_L5L6_number;
wire [9:0] FM_L5L6_L3_FromPlus_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L3_FromPlus_FT_L5L6;
wire FM_L5L6_L3_FromPlus_FT_L5L6_read_en;
FullMatch #(128) FM_L5L6_L3_FromPlus(
.data_in(MT_L5L6_Plus_FM_L5L6_L3_FromPlus),
.enable(MT_L5L6_Plus_FM_L5L6_L3_FromPlus_wr_en),
.number_out(FM_L5L6_L3_FromPlus_FT_L5L6_number),
.read_add(FM_L5L6_L3_FromPlus_FT_L5L6_read_add),
.data_out(FM_L5L6_L3_FromPlus_FT_L5L6),
.read_en(FM_L5L6_L3_FromPlus_FT_L5L6_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L5L6_Plus_FM_L5L6_L4_FromPlus;
wire MT_L5L6_Plus_FM_L5L6_L4_FromPlus_wr_en;
wire [5:0] FM_L5L6_L4_FromPlus_FT_L5L6_number;
wire [9:0] FM_L5L6_L4_FromPlus_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L4_FromPlus_FT_L5L6;
wire FM_L5L6_L4_FromPlus_FT_L5L6_read_en;
FullMatch #(128) FM_L5L6_L4_FromPlus(
.data_in(MT_L5L6_Plus_FM_L5L6_L4_FromPlus),
.enable(MT_L5L6_Plus_FM_L5L6_L4_FromPlus_wr_en),
.number_out(FM_L5L6_L4_FromPlus_FT_L5L6_number),
.read_add(FM_L5L6_L4_FromPlus_FT_L5L6_read_add),
.data_out(FM_L5L6_L4_FromPlus_FT_L5L6),
.read_en(FM_L5L6_L4_FromPlus_FT_L5L6_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L5L6_Minus_FM_L5L6_L1_FromMinus;
wire MT_L5L6_Minus_FM_L5L6_L1_FromMinus_wr_en;
wire [5:0] FM_L5L6_L1_FromMinus_FT_L5L6_number;
wire [9:0] FM_L5L6_L1_FromMinus_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L1_FromMinus_FT_L5L6;
wire FM_L5L6_L1_FromMinus_FT_L5L6_read_en;
FullMatch #(128) FM_L5L6_L1_FromMinus(
.data_in(MT_L5L6_Minus_FM_L5L6_L1_FromMinus),
.enable(MT_L5L6_Minus_FM_L5L6_L1_FromMinus_wr_en),
.number_out(FM_L5L6_L1_FromMinus_FT_L5L6_number),
.read_add(FM_L5L6_L1_FromMinus_FT_L5L6_read_add),
.data_out(FM_L5L6_L1_FromMinus_FT_L5L6),
.read_en(FM_L5L6_L1_FromMinus_FT_L5L6_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L5L6_Minus_FM_L5L6_L2_FromMinus;
wire MT_L5L6_Minus_FM_L5L6_L2_FromMinus_wr_en;
wire [5:0] FM_L5L6_L2_FromMinus_FT_L5L6_number;
wire [9:0] FM_L5L6_L2_FromMinus_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L2_FromMinus_FT_L5L6;
wire FM_L5L6_L2_FromMinus_FT_L5L6_read_en;
FullMatch #(128) FM_L5L6_L2_FromMinus(
.data_in(MT_L5L6_Minus_FM_L5L6_L2_FromMinus),
.enable(MT_L5L6_Minus_FM_L5L6_L2_FromMinus_wr_en),
.number_out(FM_L5L6_L2_FromMinus_FT_L5L6_number),
.read_add(FM_L5L6_L2_FromMinus_FT_L5L6_read_add),
.data_out(FM_L5L6_L2_FromMinus_FT_L5L6),
.read_en(FM_L5L6_L2_FromMinus_FT_L5L6_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L5L6_Minus_FM_L5L6_L3_FromMinus;
wire MT_L5L6_Minus_FM_L5L6_L3_FromMinus_wr_en;
wire [5:0] FM_L5L6_L3_FromMinus_FT_L5L6_number;
wire [9:0] FM_L5L6_L3_FromMinus_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L3_FromMinus_FT_L5L6;
wire FM_L5L6_L3_FromMinus_FT_L5L6_read_en;
FullMatch #(128) FM_L5L6_L3_FromMinus(
.data_in(MT_L5L6_Minus_FM_L5L6_L3_FromMinus),
.enable(MT_L5L6_Minus_FM_L5L6_L3_FromMinus_wr_en),
.number_out(FM_L5L6_L3_FromMinus_FT_L5L6_number),
.read_add(FM_L5L6_L3_FromMinus_FT_L5L6_read_add),
.data_out(FM_L5L6_L3_FromMinus_FT_L5L6),
.read_en(FM_L5L6_L3_FromMinus_FT_L5L6_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [35:0] MT_L5L6_Minus_FM_L5L6_L4_FromMinus;
wire MT_L5L6_Minus_FM_L5L6_L4_FromMinus_wr_en;
wire [5:0] FM_L5L6_L4_FromMinus_FT_L5L6_number;
wire [9:0] FM_L5L6_L4_FromMinus_FT_L5L6_read_add;
wire [35:0] FM_L5L6_L4_FromMinus_FT_L5L6;
wire FM_L5L6_L4_FromMinus_FT_L5L6_read_en;
FullMatch #(128) FM_L5L6_L4_FromMinus(
.data_in(MT_L5L6_Minus_FM_L5L6_L4_FromMinus),
.enable(MT_L5L6_Minus_FM_L5L6_L4_FromMinus_wr_en),
.number_out(FM_L5L6_L4_FromMinus_FT_L5L6_number),
.read_add(FM_L5L6_L4_FromMinus_FT_L5L6_read_add),
.data_out(FM_L5L6_L4_FromMinus_FT_L5L6),
.read_en(FM_L5L6_L4_FromMinus_FT_L5L6_read_en),
.start(start10_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [125:0] FT_L1L2_TF_L1L2;
wire FT_L1L2_TF_L1L2_wr_en;
//wire TF_L1L2_DataStream;
TrackFit  TF_L1L2(
.data_in(FT_L1L2_TF_L1L2),
.enable(FT_L1L2_TF_L1L2_wr_en),
.data_out(TF_L1L2_DataStream),
.start(start11_0),
.done(done10_5),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [125:0] FT_L3L4_TF_L3L4;
wire FT_L3L4_TF_L3L4_wr_en;
//wire TF_L3L4_DataStream;
TrackFit  TF_L3L4(
.data_in(FT_L3L4_TF_L3L4),
.enable(FT_L3L4_TF_L3L4_wr_en),
.data_out(TF_L3L4_DataStream),
.start(start11_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


wire [125:0] FT_L5L6_TF_L5L6;
wire FT_L5L6_TF_L5L6_wr_en;
//wire TF_L5L6_DataStream;
TrackFit  TF_L5L6(
.data_in(FT_L5L6_TF_L5L6),
.enable(FT_L5L6_TF_L5L6_wr_en),
.data_out(TF_L5L6_DataStream),
.start(start11_0),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


LayerRouter  LR1_D3(
.stubin(IL1_D3_LR1_D3),
.stuboutL1(LR1_D3_SL1_L1D3),
.stuboutL3(LR1_D3_SL1_L3D3),
.stuboutL5(LR1_D3_SL1_L5D3),
.stuboutL2(LR1_D3_SL1_L2D3),
.stuboutL4(LR1_D3_SL1_L4D3),
.stuboutL6(LR1_D3_SL1_L6D3),
.wr_en1(LR1_D3_SL1_L1D3_wr_en),
.wr_en2(LR1_D3_SL1_L3D3_wr_en),
.wr_en3(LR1_D3_SL1_L5D3_wr_en),
.wr_en4(LR1_D3_SL1_L2D3_wr_en),
.wr_en5(LR1_D3_SL1_L4D3_wr_en),
.wr_en6(LR1_D3_SL1_L6D3_wr_en),
.start(start1_5),
.done(done1_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


LayerRouter  LR2_D3(
.stubin(IL2_D3_LR2_D3),
.stuboutL1(LR2_D3_SL2_L1D3),
.stuboutL3(LR2_D3_SL2_L3D3),
.stuboutL5(LR2_D3_SL2_L5D3),
.stuboutL2(LR2_D3_SL2_L2D3),
.stuboutL4(LR2_D3_SL2_L4D3),
.stuboutL6(LR2_D3_SL2_L6D3),
.wr_en1(LR2_D3_SL2_L1D3_wr_en),
.wr_en2(LR2_D3_SL2_L3D3_wr_en),
.wr_en3(LR2_D3_SL2_L5D3_wr_en),
.wr_en4(LR2_D3_SL2_L2D3_wr_en),
.wr_en5(LR2_D3_SL2_L4D3_wr_en),
.wr_en6(LR2_D3_SL2_L6D3_wr_en),
.start(start1_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


LayerRouter  LR3_D3(
.stubin(IL3_D3_LR3_D3),
.stuboutL1(LR3_D3_SL3_L1D3),
.stuboutL3(LR3_D3_SL3_L3D3),
.stuboutL5(LR3_D3_SL3_L5D3),
.stuboutL2(LR3_D3_SL3_L2D3),
.stuboutL4(LR3_D3_SL3_L4D3),
.stuboutL6(LR3_D3_SL3_L6D3),
.wr_en1(LR3_D3_SL3_L1D3_wr_en),
.wr_en2(LR3_D3_SL3_L3D3_wr_en),
.wr_en3(LR3_D3_SL3_L5D3_wr_en),
.wr_en4(LR3_D3_SL3_L2D3_wr_en),
.wr_en5(LR3_D3_SL3_L4D3_wr_en),
.wr_en6(LR3_D3_SL3_L6D3_wr_en),
.start(start1_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


LayerRouter  LR1_D4(
.stubin(IL1_D4_LR1_D4),
.stuboutL1(LR1_D4_SL1_L1D4),
.stuboutL3(LR1_D4_SL1_L3D4),
.stuboutL5(LR1_D4_SL1_L5D4),
.stuboutL2(LR1_D4_SL1_L2D4),
.stuboutL4(LR1_D4_SL1_L4D4),
.stuboutL6(LR1_D4_SL1_L6D4),
.wr_en1(LR1_D4_SL1_L1D4_wr_en),
.wr_en2(LR1_D4_SL1_L3D4_wr_en),
.wr_en3(LR1_D4_SL1_L5D4_wr_en),
.wr_en4(LR1_D4_SL1_L2D4_wr_en),
.wr_en5(LR1_D4_SL1_L4D4_wr_en),
.wr_en6(LR1_D4_SL1_L6D4_wr_en),
.start(start1_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


LayerRouter  LR2_D4(
.stubin(IL2_D4_LR2_D4),
.stuboutL1(LR2_D4_SL2_L1D4),
.stuboutL3(LR2_D4_SL2_L3D4),
.stuboutL5(LR2_D4_SL2_L5D4),
.stuboutL2(LR2_D4_SL2_L2D4),
.stuboutL4(LR2_D4_SL2_L4D4),
.stuboutL6(LR2_D4_SL2_L6D4),
.wr_en1(LR2_D4_SL2_L1D4_wr_en),
.wr_en2(LR2_D4_SL2_L3D4_wr_en),
.wr_en3(LR2_D4_SL2_L5D4_wr_en),
.wr_en4(LR2_D4_SL2_L2D4_wr_en),
.wr_en5(LR2_D4_SL2_L4D4_wr_en),
.wr_en6(LR2_D4_SL2_L6D4_wr_en),
.start(start1_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


LayerRouter  LR3_D4(
.stubin(IL3_D4_LR3_D4),
.stuboutL1(LR3_D4_SL3_L1D4),
.stuboutL3(LR3_D4_SL3_L3D4),
.stuboutL5(LR3_D4_SL3_L5D4),
.stuboutL2(LR3_D4_SL3_L2D4),
.stuboutL4(LR3_D4_SL3_L4D4),
.stuboutL6(LR3_D4_SL3_L6D4),
.wr_en1(LR3_D4_SL3_L1D4_wr_en),
.wr_en2(LR3_D4_SL3_L3D4_wr_en),
.wr_en3(LR3_D4_SL3_L5D4_wr_en),
.wr_en4(LR3_D4_SL3_L2D4_wr_en),
.wr_en5(LR3_D4_SL3_L4D4_wr_en),
.wr_en6(LR3_D4_SL3_L6D4_wr_en),
.start(start1_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b1,1'b1) VMR_L1D3(
.number_in1(SL1_L1D3_VMR_L1D3_number),
.read_add1(SL1_L1D3_VMR_L1D3_read_add),
.stubinLink1(SL1_L1D3_VMR_L1D3),
.number_in2(SL2_L1D3_VMR_L1D3_number),
.read_add2(SL2_L1D3_VMR_L1D3_read_add),
.stubinLink2(SL2_L1D3_VMR_L1D3),
.number_in3(SL3_L1D3_VMR_L1D3_number),
.read_add3(SL3_L1D3_VMR_L1D3_read_add),
.stubinLink3(SL3_L1D3_VMR_L1D3),
.vmstuboutPHI1Z1n1(VMR_L1D3_VMS_L1D3PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L1D3_VMS_L1D3PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L1D3_VMS_L1D3PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L1D3_VMS_L1D3PHI1Z1n4),
.vmstuboutPHI1Z1n5(VMR_L1D3_VMS_L1D3PHI1Z1n5),
.vmstuboutPHI1Z1n6(VMR_L1D3_VMS_L1D3PHI1Z1n6),
.vmstuboutPHI1Z1n7(VMR_L1D3_VMS_L1D3PHI1Z1n7),
.vmstuboutPHI1Z1n8(VMR_L1D3_VMS_L1D3PHI1Z1n8),
.vmstuboutPHI2Z1n1(VMR_L1D3_VMS_L1D3PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L1D3_VMS_L1D3PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L1D3_VMS_L1D3PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L1D3_VMS_L1D3PHI2Z1n4),
.vmstuboutPHI2Z1n5(VMR_L1D3_VMS_L1D3PHI2Z1n5),
.vmstuboutPHI2Z1n6(VMR_L1D3_VMS_L1D3PHI2Z1n6),
.vmstuboutPHI2Z1n7(VMR_L1D3_VMS_L1D3PHI2Z1n7),
.vmstuboutPHI2Z1n8(VMR_L1D3_VMS_L1D3PHI2Z1n8),
.vmstuboutPHI3Z1n1(VMR_L1D3_VMS_L1D3PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L1D3_VMS_L1D3PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L1D3_VMS_L1D3PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L1D3_VMS_L1D3PHI3Z1n4),
.vmstuboutPHI3Z1n5(VMR_L1D3_VMS_L1D3PHI3Z1n5),
.vmstuboutPHI3Z1n6(VMR_L1D3_VMS_L1D3PHI3Z1n6),
.vmstuboutPHI3Z1n7(VMR_L1D3_VMS_L1D3PHI3Z1n7),
.vmstuboutPHI3Z1n8(VMR_L1D3_VMS_L1D3PHI3Z1n8),
.vmstuboutPHI1Z2n1(VMR_L1D3_VMS_L1D3PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L1D3_VMS_L1D3PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L1D3_VMS_L1D3PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L1D3_VMS_L1D3PHI1Z2n4),
.vmstuboutPHI1Z2n5(VMR_L1D3_VMS_L1D3PHI1Z2n5),
.vmstuboutPHI1Z2n6(VMR_L1D3_VMS_L1D3PHI1Z2n6),
.vmstuboutPHI1Z2n7(VMR_L1D3_VMS_L1D3PHI1Z2n7),
.vmstuboutPHI1Z2n8(VMR_L1D3_VMS_L1D3PHI1Z2n8),
.vmstuboutPHI2Z2n1(VMR_L1D3_VMS_L1D3PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L1D3_VMS_L1D3PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L1D3_VMS_L1D3PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L1D3_VMS_L1D3PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L1D3_VMS_L1D3PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L1D3_VMS_L1D3PHI2Z2n6),
.vmstuboutPHI2Z2n7(VMR_L1D3_VMS_L1D3PHI2Z2n7),
.vmstuboutPHI2Z2n8(VMR_L1D3_VMS_L1D3PHI2Z2n8),
.vmstuboutPHI3Z2n1(VMR_L1D3_VMS_L1D3PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L1D3_VMS_L1D3PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L1D3_VMS_L1D3PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L1D3_VMS_L1D3PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L1D3_VMS_L1D3PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L1D3_VMS_L1D3PHI3Z2n6),
.vmstuboutPHI3Z2n7(VMR_L1D3_VMS_L1D3PHI3Z2n7),
.vmstuboutPHI3Z2n8(VMR_L1D3_VMS_L1D3PHI3Z2n8),
.allstuboutn1(VMR_L1D3_AS_L1D3n1),
.allstuboutn2(VMR_L1D3_AS_L1D3n2),
.allstuboutn3(VMR_L1D3_AS_L1D3n3),
.allstuboutn4(VMR_L1D3_AS_L1D3n4),
.vmstuboutPHI1Z1n1_wr_en(VMR_L1D3_VMS_L1D3PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L1D3_VMS_L1D3PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L1D3_VMS_L1D3PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L1D3_VMS_L1D3PHI1Z1n4_wr_en),
.vmstuboutPHI1Z1n5_wr_en(VMR_L1D3_VMS_L1D3PHI1Z1n5_wr_en),
.vmstuboutPHI1Z1n6_wr_en(VMR_L1D3_VMS_L1D3PHI1Z1n6_wr_en),
.vmstuboutPHI1Z1n7_wr_en(VMR_L1D3_VMS_L1D3PHI1Z1n7_wr_en),
.vmstuboutPHI1Z1n8_wr_en(VMR_L1D3_VMS_L1D3PHI1Z1n8_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L1D3_VMS_L1D3PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L1D3_VMS_L1D3PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L1D3_VMS_L1D3PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L1D3_VMS_L1D3PHI2Z1n4_wr_en),
.vmstuboutPHI2Z1n5_wr_en(VMR_L1D3_VMS_L1D3PHI2Z1n5_wr_en),
.vmstuboutPHI2Z1n6_wr_en(VMR_L1D3_VMS_L1D3PHI2Z1n6_wr_en),
.vmstuboutPHI2Z1n7_wr_en(VMR_L1D3_VMS_L1D3PHI2Z1n7_wr_en),
.vmstuboutPHI2Z1n8_wr_en(VMR_L1D3_VMS_L1D3PHI2Z1n8_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L1D3_VMS_L1D3PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L1D3_VMS_L1D3PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L1D3_VMS_L1D3PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L1D3_VMS_L1D3PHI3Z1n4_wr_en),
.vmstuboutPHI3Z1n5_wr_en(VMR_L1D3_VMS_L1D3PHI3Z1n5_wr_en),
.vmstuboutPHI3Z1n6_wr_en(VMR_L1D3_VMS_L1D3PHI3Z1n6_wr_en),
.vmstuboutPHI3Z1n7_wr_en(VMR_L1D3_VMS_L1D3PHI3Z1n7_wr_en),
.vmstuboutPHI3Z1n8_wr_en(VMR_L1D3_VMS_L1D3PHI3Z1n8_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L1D3_VMS_L1D3PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L1D3_VMS_L1D3PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L1D3_VMS_L1D3PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L1D3_VMS_L1D3PHI1Z2n4_wr_en),
.vmstuboutPHI1Z2n5_wr_en(VMR_L1D3_VMS_L1D3PHI1Z2n5_wr_en),
.vmstuboutPHI1Z2n6_wr_en(VMR_L1D3_VMS_L1D3PHI1Z2n6_wr_en),
.vmstuboutPHI1Z2n7_wr_en(VMR_L1D3_VMS_L1D3PHI1Z2n7_wr_en),
.vmstuboutPHI1Z2n8_wr_en(VMR_L1D3_VMS_L1D3PHI1Z2n8_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L1D3_VMS_L1D3PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L1D3_VMS_L1D3PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L1D3_VMS_L1D3PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L1D3_VMS_L1D3PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L1D3_VMS_L1D3PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L1D3_VMS_L1D3PHI2Z2n6_wr_en),
.vmstuboutPHI2Z2n7_wr_en(VMR_L1D3_VMS_L1D3PHI2Z2n7_wr_en),
.vmstuboutPHI2Z2n8_wr_en(VMR_L1D3_VMS_L1D3PHI2Z2n8_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L1D3_VMS_L1D3PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L1D3_VMS_L1D3PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L1D3_VMS_L1D3PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L1D3_VMS_L1D3PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L1D3_VMS_L1D3PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L1D3_VMS_L1D3PHI3Z2n6_wr_en),
.vmstuboutPHI3Z2n7_wr_en(VMR_L1D3_VMS_L1D3PHI3Z2n7_wr_en),
.vmstuboutPHI3Z2n8_wr_en(VMR_L1D3_VMS_L1D3PHI3Z2n8_wr_en),
.valid_data1(VMR_L1D3_AS_L1D3n1_wr_en),
.valid_data2(VMR_L1D3_AS_L1D3n2_wr_en),
.valid_data3(VMR_L1D3_AS_L1D3n3_wr_en),
.valid_data4(VMR_L1D3_AS_L1D3n4_wr_en),
.start(start2_5),
.done(done2_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b1,1'b1) VMR_L1D4(
.number_in1(SL1_L1D4_VMR_L1D4_number),
.read_add1(SL1_L1D4_VMR_L1D4_read_add),
.stubinLink1(SL1_L1D4_VMR_L1D4),
.number_in2(SL2_L1D4_VMR_L1D4_number),
.read_add2(SL2_L1D4_VMR_L1D4_read_add),
.stubinLink2(SL2_L1D4_VMR_L1D4),
.number_in3(SL3_L1D4_VMR_L1D4_number),
.read_add3(SL3_L1D4_VMR_L1D4_read_add),
.stubinLink3(SL3_L1D4_VMR_L1D4),
.vmstuboutPHI1Z1n1(VMR_L1D4_VMS_L1D4PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L1D4_VMS_L1D4PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L1D4_VMS_L1D4PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L1D4_VMS_L1D4PHI1Z1n4),
.vmstuboutPHI2Z1n1(VMR_L1D4_VMS_L1D4PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L1D4_VMS_L1D4PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L1D4_VMS_L1D4PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L1D4_VMS_L1D4PHI2Z1n4),
.vmstuboutPHI3Z1n1(VMR_L1D4_VMS_L1D4PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L1D4_VMS_L1D4PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L1D4_VMS_L1D4PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L1D4_VMS_L1D4PHI3Z1n4),
.allstuboutn1(VMR_L1D4_AS_L1D4n1),
.allstuboutn2(VMR_L1D4_AS_L1D4n2),
.allstuboutn3(VMR_L1D4_AS_L1D4n3),
.vmstuboutPHI1Z2n1(VMR_L1D4_VMS_L1D4PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L1D4_VMS_L1D4PHI1Z2n2),
.vmstuboutPHI2Z2n1(VMR_L1D4_VMS_L1D4PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L1D4_VMS_L1D4PHI2Z2n2),
.vmstuboutPHI3Z2n1(VMR_L1D4_VMS_L1D4PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L1D4_VMS_L1D4PHI3Z2n2),
.vmstuboutPHI1Z1n1_wr_en(VMR_L1D4_VMS_L1D4PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L1D4_VMS_L1D4PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L1D4_VMS_L1D4PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L1D4_VMS_L1D4PHI1Z1n4_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L1D4_VMS_L1D4PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L1D4_VMS_L1D4PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L1D4_VMS_L1D4PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L1D4_VMS_L1D4PHI2Z1n4_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L1D4_VMS_L1D4PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L1D4_VMS_L1D4PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L1D4_VMS_L1D4PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L1D4_VMS_L1D4PHI3Z1n4_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L1D4_VMS_L1D4PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L1D4_VMS_L1D4PHI1Z2n2_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L1D4_VMS_L1D4PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L1D4_VMS_L1D4PHI2Z2n2_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L1D4_VMS_L1D4PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L1D4_VMS_L1D4PHI3Z2n2_wr_en),
.valid_data1(VMR_L1D4_AS_L1D4n1_wr_en),
.valid_data2(VMR_L1D4_AS_L1D4n2_wr_en),
.valid_data3(VMR_L1D4_AS_L1D4n3_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b1,1'b1) VMR_L3D3(
.number_in1(SL1_L3D3_VMR_L3D3_number),
.read_add1(SL1_L3D3_VMR_L3D3_read_add),
.stubinLink1(SL1_L3D3_VMR_L3D3),
.number_in2(SL2_L3D3_VMR_L3D3_number),
.read_add2(SL2_L3D3_VMR_L3D3_read_add),
.stubinLink2(SL2_L3D3_VMR_L3D3),
.number_in3(SL3_L3D3_VMR_L3D3_number),
.read_add3(SL3_L3D3_VMR_L3D3_read_add),
.stubinLink3(SL3_L3D3_VMR_L3D3),
.vmstuboutPHI1Z1n1(VMR_L3D3_VMS_L3D3PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L3D3_VMS_L3D3PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L3D3_VMS_L3D3PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L3D3_VMS_L3D3PHI1Z1n4),
.vmstuboutPHI1Z1n5(VMR_L3D3_VMS_L3D3PHI1Z1n5),
.vmstuboutPHI1Z1n6(VMR_L3D3_VMS_L3D3PHI1Z1n6),
.vmstuboutPHI2Z1n1(VMR_L3D3_VMS_L3D3PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L3D3_VMS_L3D3PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L3D3_VMS_L3D3PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L3D3_VMS_L3D3PHI2Z1n4),
.vmstuboutPHI2Z1n5(VMR_L3D3_VMS_L3D3PHI2Z1n5),
.vmstuboutPHI2Z1n6(VMR_L3D3_VMS_L3D3PHI2Z1n6),
.vmstuboutPHI3Z1n1(VMR_L3D3_VMS_L3D3PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L3D3_VMS_L3D3PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L3D3_VMS_L3D3PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L3D3_VMS_L3D3PHI3Z1n4),
.vmstuboutPHI3Z1n5(VMR_L3D3_VMS_L3D3PHI3Z1n5),
.vmstuboutPHI3Z1n6(VMR_L3D3_VMS_L3D3PHI3Z1n6),
.vmstuboutPHI1Z2n1(VMR_L3D3_VMS_L3D3PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L3D3_VMS_L3D3PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L3D3_VMS_L3D3PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L3D3_VMS_L3D3PHI1Z2n4),
.vmstuboutPHI1Z2n5(VMR_L3D3_VMS_L3D3PHI1Z2n5),
.vmstuboutPHI1Z2n6(VMR_L3D3_VMS_L3D3PHI1Z2n6),
.vmstuboutPHI2Z2n1(VMR_L3D3_VMS_L3D3PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L3D3_VMS_L3D3PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L3D3_VMS_L3D3PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L3D3_VMS_L3D3PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L3D3_VMS_L3D3PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L3D3_VMS_L3D3PHI2Z2n6),
.vmstuboutPHI3Z2n1(VMR_L3D3_VMS_L3D3PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L3D3_VMS_L3D3PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L3D3_VMS_L3D3PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L3D3_VMS_L3D3PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L3D3_VMS_L3D3PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L3D3_VMS_L3D3PHI3Z2n6),
.allstuboutn1(VMR_L3D3_AS_L3D3n1),
.allstuboutn2(VMR_L3D3_AS_L3D3n2),
.allstuboutn3(VMR_L3D3_AS_L3D3n3),
.allstuboutn4(VMR_L3D3_AS_L3D3n4),
.vmstuboutPHI1Z1n1_wr_en(VMR_L3D3_VMS_L3D3PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L3D3_VMS_L3D3PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L3D3_VMS_L3D3PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L3D3_VMS_L3D3PHI1Z1n4_wr_en),
.vmstuboutPHI1Z1n5_wr_en(VMR_L3D3_VMS_L3D3PHI1Z1n5_wr_en),
.vmstuboutPHI1Z1n6_wr_en(VMR_L3D3_VMS_L3D3PHI1Z1n6_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L3D3_VMS_L3D3PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L3D3_VMS_L3D3PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L3D3_VMS_L3D3PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L3D3_VMS_L3D3PHI2Z1n4_wr_en),
.vmstuboutPHI2Z1n5_wr_en(VMR_L3D3_VMS_L3D3PHI2Z1n5_wr_en),
.vmstuboutPHI2Z1n6_wr_en(VMR_L3D3_VMS_L3D3PHI2Z1n6_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L3D3_VMS_L3D3PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L3D3_VMS_L3D3PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L3D3_VMS_L3D3PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L3D3_VMS_L3D3PHI3Z1n4_wr_en),
.vmstuboutPHI3Z1n5_wr_en(VMR_L3D3_VMS_L3D3PHI3Z1n5_wr_en),
.vmstuboutPHI3Z1n6_wr_en(VMR_L3D3_VMS_L3D3PHI3Z1n6_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L3D3_VMS_L3D3PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L3D3_VMS_L3D3PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L3D3_VMS_L3D3PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L3D3_VMS_L3D3PHI1Z2n4_wr_en),
.vmstuboutPHI1Z2n5_wr_en(VMR_L3D3_VMS_L3D3PHI1Z2n5_wr_en),
.vmstuboutPHI1Z2n6_wr_en(VMR_L3D3_VMS_L3D3PHI1Z2n6_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L3D3_VMS_L3D3PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L3D3_VMS_L3D3PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L3D3_VMS_L3D3PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L3D3_VMS_L3D3PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L3D3_VMS_L3D3PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L3D3_VMS_L3D3PHI2Z2n6_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L3D3_VMS_L3D3PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L3D3_VMS_L3D3PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L3D3_VMS_L3D3PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L3D3_VMS_L3D3PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L3D3_VMS_L3D3PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L3D3_VMS_L3D3PHI3Z2n6_wr_en),
.valid_data1(VMR_L3D3_AS_L3D3n1_wr_en),
.valid_data2(VMR_L3D3_AS_L3D3n2_wr_en),
.valid_data3(VMR_L3D3_AS_L3D3n3_wr_en),
.valid_data4(VMR_L3D3_AS_L3D3n4_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b1,1'b1) VMR_L3D4(
.number_in1(SL1_L3D4_VMR_L3D4_number),
.read_add1(SL1_L3D4_VMR_L3D4_read_add),
.stubinLink1(SL1_L3D4_VMR_L3D4),
.number_in2(SL2_L3D4_VMR_L3D4_number),
.read_add2(SL2_L3D4_VMR_L3D4_read_add),
.stubinLink2(SL2_L3D4_VMR_L3D4),
.number_in3(SL3_L3D4_VMR_L3D4_number),
.read_add3(SL3_L3D4_VMR_L3D4_read_add),
.stubinLink3(SL3_L3D4_VMR_L3D4),
.vmstuboutPHI1Z1n1(VMR_L3D4_VMS_L3D4PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L3D4_VMS_L3D4PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L3D4_VMS_L3D4PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L3D4_VMS_L3D4PHI1Z1n4),
.vmstuboutPHI1Z1n5(VMR_L3D4_VMS_L3D4PHI1Z1n5),
.vmstuboutPHI1Z1n6(VMR_L3D4_VMS_L3D4PHI1Z1n6),
.vmstuboutPHI2Z1n1(VMR_L3D4_VMS_L3D4PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L3D4_VMS_L3D4PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L3D4_VMS_L3D4PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L3D4_VMS_L3D4PHI2Z1n4),
.vmstuboutPHI2Z1n5(VMR_L3D4_VMS_L3D4PHI2Z1n5),
.vmstuboutPHI2Z1n6(VMR_L3D4_VMS_L3D4PHI2Z1n6),
.vmstuboutPHI3Z1n1(VMR_L3D4_VMS_L3D4PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L3D4_VMS_L3D4PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L3D4_VMS_L3D4PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L3D4_VMS_L3D4PHI3Z1n4),
.vmstuboutPHI3Z1n5(VMR_L3D4_VMS_L3D4PHI3Z1n5),
.vmstuboutPHI3Z1n6(VMR_L3D4_VMS_L3D4PHI3Z1n6),
.vmstuboutPHI1Z2n1(VMR_L3D4_VMS_L3D4PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L3D4_VMS_L3D4PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L3D4_VMS_L3D4PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L3D4_VMS_L3D4PHI1Z2n4),
.vmstuboutPHI2Z2n1(VMR_L3D4_VMS_L3D4PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L3D4_VMS_L3D4PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L3D4_VMS_L3D4PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L3D4_VMS_L3D4PHI2Z2n4),
.vmstuboutPHI3Z2n1(VMR_L3D4_VMS_L3D4PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L3D4_VMS_L3D4PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L3D4_VMS_L3D4PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L3D4_VMS_L3D4PHI3Z2n4),
.allstuboutn1(VMR_L3D4_AS_L3D4n1),
.allstuboutn2(VMR_L3D4_AS_L3D4n2),
.allstuboutn3(VMR_L3D4_AS_L3D4n3),
.vmstuboutPHI1Z1n1_wr_en(VMR_L3D4_VMS_L3D4PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L3D4_VMS_L3D4PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L3D4_VMS_L3D4PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L3D4_VMS_L3D4PHI1Z1n4_wr_en),
.vmstuboutPHI1Z1n5_wr_en(VMR_L3D4_VMS_L3D4PHI1Z1n5_wr_en),
.vmstuboutPHI1Z1n6_wr_en(VMR_L3D4_VMS_L3D4PHI1Z1n6_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L3D4_VMS_L3D4PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L3D4_VMS_L3D4PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L3D4_VMS_L3D4PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L3D4_VMS_L3D4PHI2Z1n4_wr_en),
.vmstuboutPHI2Z1n5_wr_en(VMR_L3D4_VMS_L3D4PHI2Z1n5_wr_en),
.vmstuboutPHI2Z1n6_wr_en(VMR_L3D4_VMS_L3D4PHI2Z1n6_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L3D4_VMS_L3D4PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L3D4_VMS_L3D4PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L3D4_VMS_L3D4PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L3D4_VMS_L3D4PHI3Z1n4_wr_en),
.vmstuboutPHI3Z1n5_wr_en(VMR_L3D4_VMS_L3D4PHI3Z1n5_wr_en),
.vmstuboutPHI3Z1n6_wr_en(VMR_L3D4_VMS_L3D4PHI3Z1n6_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L3D4_VMS_L3D4PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L3D4_VMS_L3D4PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L3D4_VMS_L3D4PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L3D4_VMS_L3D4PHI1Z2n4_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L3D4_VMS_L3D4PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L3D4_VMS_L3D4PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L3D4_VMS_L3D4PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L3D4_VMS_L3D4PHI2Z2n4_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L3D4_VMS_L3D4PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L3D4_VMS_L3D4PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L3D4_VMS_L3D4PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L3D4_VMS_L3D4PHI3Z2n4_wr_en),
.valid_data1(VMR_L3D4_AS_L3D4n1_wr_en),
.valid_data2(VMR_L3D4_AS_L3D4n2_wr_en),
.valid_data3(VMR_L3D4_AS_L3D4n3_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b0,1'b1) VMR_L5D3(
.number_in1(SL1_L5D3_VMR_L5D3_number),
.read_add1(SL1_L5D3_VMR_L5D3_read_add),
.stubinLink1(SL1_L5D3_VMR_L5D3),
.number_in2(SL2_L5D3_VMR_L5D3_number),
.read_add2(SL2_L5D3_VMR_L5D3_read_add),
.stubinLink2(SL2_L5D3_VMR_L5D3),
.number_in3(SL3_L5D3_VMR_L5D3_number),
.read_add3(SL3_L5D3_VMR_L5D3_read_add),
.stubinLink3(SL3_L5D3_VMR_L5D3),
.vmstuboutPHI1Z1n1(VMR_L5D3_VMS_L5D3PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L5D3_VMS_L5D3PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L5D3_VMS_L5D3PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L5D3_VMS_L5D3PHI1Z1n4),
.vmstuboutPHI1Z1n5(VMR_L5D3_VMS_L5D3PHI1Z1n5),
.vmstuboutPHI1Z1n6(VMR_L5D3_VMS_L5D3PHI1Z1n6),
.vmstuboutPHI2Z1n1(VMR_L5D3_VMS_L5D3PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L5D3_VMS_L5D3PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L5D3_VMS_L5D3PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L5D3_VMS_L5D3PHI2Z1n4),
.vmstuboutPHI2Z1n5(VMR_L5D3_VMS_L5D3PHI2Z1n5),
.vmstuboutPHI2Z1n6(VMR_L5D3_VMS_L5D3PHI2Z1n6),
.vmstuboutPHI3Z1n1(VMR_L5D3_VMS_L5D3PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L5D3_VMS_L5D3PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L5D3_VMS_L5D3PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L5D3_VMS_L5D3PHI3Z1n4),
.vmstuboutPHI3Z1n5(VMR_L5D3_VMS_L5D3PHI3Z1n5),
.vmstuboutPHI3Z1n6(VMR_L5D3_VMS_L5D3PHI3Z1n6),
.vmstuboutPHI1Z2n1(VMR_L5D3_VMS_L5D3PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L5D3_VMS_L5D3PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L5D3_VMS_L5D3PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L5D3_VMS_L5D3PHI1Z2n4),
.vmstuboutPHI1Z2n5(VMR_L5D3_VMS_L5D3PHI1Z2n5),
.vmstuboutPHI1Z2n6(VMR_L5D3_VMS_L5D3PHI1Z2n6),
.vmstuboutPHI2Z2n1(VMR_L5D3_VMS_L5D3PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L5D3_VMS_L5D3PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L5D3_VMS_L5D3PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L5D3_VMS_L5D3PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L5D3_VMS_L5D3PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L5D3_VMS_L5D3PHI2Z2n6),
.vmstuboutPHI3Z2n1(VMR_L5D3_VMS_L5D3PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L5D3_VMS_L5D3PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L5D3_VMS_L5D3PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L5D3_VMS_L5D3PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L5D3_VMS_L5D3PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L5D3_VMS_L5D3PHI3Z2n6),
.allstuboutn1(VMR_L5D3_AS_L5D3n1),
.allstuboutn2(VMR_L5D3_AS_L5D3n2),
.allstuboutn3(VMR_L5D3_AS_L5D3n3),
.allstuboutn4(VMR_L5D3_AS_L5D3n4),
.vmstuboutPHI1Z1n1_wr_en(VMR_L5D3_VMS_L5D3PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L5D3_VMS_L5D3PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L5D3_VMS_L5D3PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L5D3_VMS_L5D3PHI1Z1n4_wr_en),
.vmstuboutPHI1Z1n5_wr_en(VMR_L5D3_VMS_L5D3PHI1Z1n5_wr_en),
.vmstuboutPHI1Z1n6_wr_en(VMR_L5D3_VMS_L5D3PHI1Z1n6_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L5D3_VMS_L5D3PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L5D3_VMS_L5D3PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L5D3_VMS_L5D3PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L5D3_VMS_L5D3PHI2Z1n4_wr_en),
.vmstuboutPHI2Z1n5_wr_en(VMR_L5D3_VMS_L5D3PHI2Z1n5_wr_en),
.vmstuboutPHI2Z1n6_wr_en(VMR_L5D3_VMS_L5D3PHI2Z1n6_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L5D3_VMS_L5D3PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L5D3_VMS_L5D3PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L5D3_VMS_L5D3PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L5D3_VMS_L5D3PHI3Z1n4_wr_en),
.vmstuboutPHI3Z1n5_wr_en(VMR_L5D3_VMS_L5D3PHI3Z1n5_wr_en),
.vmstuboutPHI3Z1n6_wr_en(VMR_L5D3_VMS_L5D3PHI3Z1n6_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L5D3_VMS_L5D3PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L5D3_VMS_L5D3PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L5D3_VMS_L5D3PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L5D3_VMS_L5D3PHI1Z2n4_wr_en),
.vmstuboutPHI1Z2n5_wr_en(VMR_L5D3_VMS_L5D3PHI1Z2n5_wr_en),
.vmstuboutPHI1Z2n6_wr_en(VMR_L5D3_VMS_L5D3PHI1Z2n6_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L5D3_VMS_L5D3PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L5D3_VMS_L5D3PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L5D3_VMS_L5D3PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L5D3_VMS_L5D3PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L5D3_VMS_L5D3PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L5D3_VMS_L5D3PHI2Z2n6_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L5D3_VMS_L5D3PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L5D3_VMS_L5D3PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L5D3_VMS_L5D3PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L5D3_VMS_L5D3PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L5D3_VMS_L5D3PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L5D3_VMS_L5D3PHI3Z2n6_wr_en),
.valid_data1(VMR_L5D3_AS_L5D3n1_wr_en),
.valid_data2(VMR_L5D3_AS_L5D3n2_wr_en),
.valid_data3(VMR_L5D3_AS_L5D3n3_wr_en),
.valid_data4(VMR_L5D3_AS_L5D3n4_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b0,1'b1) VMR_L5D4(
.number_in1(SL1_L5D4_VMR_L5D4_number),
.read_add1(SL1_L5D4_VMR_L5D4_read_add),
.stubinLink1(SL1_L5D4_VMR_L5D4),
.number_in2(SL2_L5D4_VMR_L5D4_number),
.read_add2(SL2_L5D4_VMR_L5D4_read_add),
.stubinLink2(SL2_L5D4_VMR_L5D4),
.number_in3(SL3_L5D4_VMR_L5D4_number),
.read_add3(SL3_L5D4_VMR_L5D4_read_add),
.stubinLink3(SL3_L5D4_VMR_L5D4),
.vmstuboutPHI1Z1n1(VMR_L5D4_VMS_L5D4PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L5D4_VMS_L5D4PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L5D4_VMS_L5D4PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L5D4_VMS_L5D4PHI1Z1n4),
.vmstuboutPHI1Z1n5(VMR_L5D4_VMS_L5D4PHI1Z1n5),
.vmstuboutPHI1Z1n6(VMR_L5D4_VMS_L5D4PHI1Z1n6),
.vmstuboutPHI2Z1n1(VMR_L5D4_VMS_L5D4PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L5D4_VMS_L5D4PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L5D4_VMS_L5D4PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L5D4_VMS_L5D4PHI2Z1n4),
.vmstuboutPHI2Z1n5(VMR_L5D4_VMS_L5D4PHI2Z1n5),
.vmstuboutPHI2Z1n6(VMR_L5D4_VMS_L5D4PHI2Z1n6),
.vmstuboutPHI3Z1n1(VMR_L5D4_VMS_L5D4PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L5D4_VMS_L5D4PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L5D4_VMS_L5D4PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L5D4_VMS_L5D4PHI3Z1n4),
.vmstuboutPHI3Z1n5(VMR_L5D4_VMS_L5D4PHI3Z1n5),
.vmstuboutPHI3Z1n6(VMR_L5D4_VMS_L5D4PHI3Z1n6),
.vmstuboutPHI1Z2n1(VMR_L5D4_VMS_L5D4PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L5D4_VMS_L5D4PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L5D4_VMS_L5D4PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L5D4_VMS_L5D4PHI1Z2n4),
.vmstuboutPHI2Z2n1(VMR_L5D4_VMS_L5D4PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L5D4_VMS_L5D4PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L5D4_VMS_L5D4PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L5D4_VMS_L5D4PHI2Z2n4),
.vmstuboutPHI3Z2n1(VMR_L5D4_VMS_L5D4PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L5D4_VMS_L5D4PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L5D4_VMS_L5D4PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L5D4_VMS_L5D4PHI3Z2n4),
.allstuboutn1(VMR_L5D4_AS_L5D4n1),
.allstuboutn2(VMR_L5D4_AS_L5D4n2),
.allstuboutn3(VMR_L5D4_AS_L5D4n3),
.vmstuboutPHI1Z1n1_wr_en(VMR_L5D4_VMS_L5D4PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L5D4_VMS_L5D4PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L5D4_VMS_L5D4PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L5D4_VMS_L5D4PHI1Z1n4_wr_en),
.vmstuboutPHI1Z1n5_wr_en(VMR_L5D4_VMS_L5D4PHI1Z1n5_wr_en),
.vmstuboutPHI1Z1n6_wr_en(VMR_L5D4_VMS_L5D4PHI1Z1n6_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L5D4_VMS_L5D4PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L5D4_VMS_L5D4PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L5D4_VMS_L5D4PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L5D4_VMS_L5D4PHI2Z1n4_wr_en),
.vmstuboutPHI2Z1n5_wr_en(VMR_L5D4_VMS_L5D4PHI2Z1n5_wr_en),
.vmstuboutPHI2Z1n6_wr_en(VMR_L5D4_VMS_L5D4PHI2Z1n6_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L5D4_VMS_L5D4PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L5D4_VMS_L5D4PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L5D4_VMS_L5D4PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L5D4_VMS_L5D4PHI3Z1n4_wr_en),
.vmstuboutPHI3Z1n5_wr_en(VMR_L5D4_VMS_L5D4PHI3Z1n5_wr_en),
.vmstuboutPHI3Z1n6_wr_en(VMR_L5D4_VMS_L5D4PHI3Z1n6_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L5D4_VMS_L5D4PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L5D4_VMS_L5D4PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L5D4_VMS_L5D4PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L5D4_VMS_L5D4PHI1Z2n4_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L5D4_VMS_L5D4PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L5D4_VMS_L5D4PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L5D4_VMS_L5D4PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L5D4_VMS_L5D4PHI2Z2n4_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L5D4_VMS_L5D4PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L5D4_VMS_L5D4PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L5D4_VMS_L5D4PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L5D4_VMS_L5D4PHI3Z2n4_wr_en),
.valid_data1(VMR_L5D4_AS_L5D4n1_wr_en),
.valid_data2(VMR_L5D4_AS_L5D4n2_wr_en),
.valid_data3(VMR_L5D4_AS_L5D4n3_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b1,1'b0) VMR_L2D3(
.number_in1(SL1_L2D3_VMR_L2D3_number),
.read_add1(SL1_L2D3_VMR_L2D3_read_add),
.stubinLink1(SL1_L2D3_VMR_L2D3),
.number_in2(SL2_L2D3_VMR_L2D3_number),
.read_add2(SL2_L2D3_VMR_L2D3_read_add),
.stubinLink2(SL2_L2D3_VMR_L2D3),
.number_in3(SL3_L2D3_VMR_L2D3_number),
.read_add3(SL3_L2D3_VMR_L2D3_read_add),
.stubinLink3(SL3_L2D3_VMR_L2D3),
.vmstuboutPHI1Z1n1(VMR_L2D3_VMS_L2D3PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L2D3_VMS_L2D3PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L2D3_VMS_L2D3PHI1Z1n3),
.vmstuboutPHI2Z1n1(VMR_L2D3_VMS_L2D3PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L2D3_VMS_L2D3PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L2D3_VMS_L2D3PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L2D3_VMS_L2D3PHI2Z1n4),
.vmstuboutPHI3Z1n1(VMR_L2D3_VMS_L2D3PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L2D3_VMS_L2D3PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L2D3_VMS_L2D3PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L2D3_VMS_L2D3PHI3Z1n4),
.vmstuboutPHI4Z1n1(VMR_L2D3_VMS_L2D3PHI4Z1n1),
.vmstuboutPHI4Z1n2(VMR_L2D3_VMS_L2D3PHI4Z1n2),
.vmstuboutPHI4Z1n3(VMR_L2D3_VMS_L2D3PHI4Z1n3),
.vmstuboutPHI1Z2n1(VMR_L2D3_VMS_L2D3PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L2D3_VMS_L2D3PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L2D3_VMS_L2D3PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L2D3_VMS_L2D3PHI1Z2n4),
.vmstuboutPHI2Z2n1(VMR_L2D3_VMS_L2D3PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L2D3_VMS_L2D3PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L2D3_VMS_L2D3PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L2D3_VMS_L2D3PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L2D3_VMS_L2D3PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L2D3_VMS_L2D3PHI2Z2n6),
.vmstuboutPHI3Z2n1(VMR_L2D3_VMS_L2D3PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L2D3_VMS_L2D3PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L2D3_VMS_L2D3PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L2D3_VMS_L2D3PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L2D3_VMS_L2D3PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L2D3_VMS_L2D3PHI3Z2n6),
.vmstuboutPHI4Z2n1(VMR_L2D3_VMS_L2D3PHI4Z2n1),
.vmstuboutPHI4Z2n2(VMR_L2D3_VMS_L2D3PHI4Z2n2),
.vmstuboutPHI4Z2n3(VMR_L2D3_VMS_L2D3PHI4Z2n3),
.vmstuboutPHI4Z2n4(VMR_L2D3_VMS_L2D3PHI4Z2n4),
.allstuboutn1(VMR_L2D3_AS_L2D3n1),
.allstuboutn2(VMR_L2D3_AS_L2D3n2),
.allstuboutn3(VMR_L2D3_AS_L2D3n3),
.vmstuboutPHI1Z1n1_wr_en(VMR_L2D3_VMS_L2D3PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L2D3_VMS_L2D3PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L2D3_VMS_L2D3PHI1Z1n3_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L2D3_VMS_L2D3PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L2D3_VMS_L2D3PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L2D3_VMS_L2D3PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L2D3_VMS_L2D3PHI2Z1n4_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L2D3_VMS_L2D3PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L2D3_VMS_L2D3PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L2D3_VMS_L2D3PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L2D3_VMS_L2D3PHI3Z1n4_wr_en),
.vmstuboutPHI4Z1n1_wr_en(VMR_L2D3_VMS_L2D3PHI4Z1n1_wr_en),
.vmstuboutPHI4Z1n2_wr_en(VMR_L2D3_VMS_L2D3PHI4Z1n2_wr_en),
.vmstuboutPHI4Z1n3_wr_en(VMR_L2D3_VMS_L2D3PHI4Z1n3_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L2D3_VMS_L2D3PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L2D3_VMS_L2D3PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L2D3_VMS_L2D3PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L2D3_VMS_L2D3PHI1Z2n4_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L2D3_VMS_L2D3PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L2D3_VMS_L2D3PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L2D3_VMS_L2D3PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L2D3_VMS_L2D3PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L2D3_VMS_L2D3PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L2D3_VMS_L2D3PHI2Z2n6_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L2D3_VMS_L2D3PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L2D3_VMS_L2D3PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L2D3_VMS_L2D3PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L2D3_VMS_L2D3PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L2D3_VMS_L2D3PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L2D3_VMS_L2D3PHI3Z2n6_wr_en),
.vmstuboutPHI4Z2n1_wr_en(VMR_L2D3_VMS_L2D3PHI4Z2n1_wr_en),
.vmstuboutPHI4Z2n2_wr_en(VMR_L2D3_VMS_L2D3PHI4Z2n2_wr_en),
.vmstuboutPHI4Z2n3_wr_en(VMR_L2D3_VMS_L2D3PHI4Z2n3_wr_en),
.vmstuboutPHI4Z2n4_wr_en(VMR_L2D3_VMS_L2D3PHI4Z2n4_wr_en),
.valid_data1(VMR_L2D3_AS_L2D3n1_wr_en),
.valid_data2(VMR_L2D3_AS_L2D3n2_wr_en),
.valid_data3(VMR_L2D3_AS_L2D3n3_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b1,1'b0) VMR_L2D4(
.number_in1(SL1_L2D4_VMR_L2D4_number),
.read_add1(SL1_L2D4_VMR_L2D4_read_add),
.stubinLink1(SL1_L2D4_VMR_L2D4),
.number_in2(SL2_L2D4_VMR_L2D4_number),
.read_add2(SL2_L2D4_VMR_L2D4_read_add),
.stubinLink2(SL2_L2D4_VMR_L2D4),
.number_in3(SL3_L2D4_VMR_L2D4_number),
.read_add3(SL3_L2D4_VMR_L2D4_read_add),
.stubinLink3(SL3_L2D4_VMR_L2D4),
.vmstuboutPHI1Z1n1(VMR_L2D4_VMS_L2D4PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L2D4_VMS_L2D4PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L2D4_VMS_L2D4PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L2D4_VMS_L2D4PHI1Z1n4),
.vmstuboutPHI2Z1n1(VMR_L2D4_VMS_L2D4PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L2D4_VMS_L2D4PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L2D4_VMS_L2D4PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L2D4_VMS_L2D4PHI2Z1n4),
.vmstuboutPHI2Z1n5(VMR_L2D4_VMS_L2D4PHI2Z1n5),
.vmstuboutPHI2Z1n6(VMR_L2D4_VMS_L2D4PHI2Z1n6),
.vmstuboutPHI3Z1n1(VMR_L2D4_VMS_L2D4PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L2D4_VMS_L2D4PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L2D4_VMS_L2D4PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L2D4_VMS_L2D4PHI3Z1n4),
.vmstuboutPHI3Z1n5(VMR_L2D4_VMS_L2D4PHI3Z1n5),
.vmstuboutPHI3Z1n6(VMR_L2D4_VMS_L2D4PHI3Z1n6),
.vmstuboutPHI4Z1n1(VMR_L2D4_VMS_L2D4PHI4Z1n1),
.vmstuboutPHI4Z1n2(VMR_L2D4_VMS_L2D4PHI4Z1n2),
.vmstuboutPHI4Z1n3(VMR_L2D4_VMS_L2D4PHI4Z1n3),
.vmstuboutPHI4Z1n4(VMR_L2D4_VMS_L2D4PHI4Z1n4),
.vmstuboutPHI1Z2n1(VMR_L2D4_VMS_L2D4PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L2D4_VMS_L2D4PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L2D4_VMS_L2D4PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L2D4_VMS_L2D4PHI1Z2n4),
.vmstuboutPHI2Z2n1(VMR_L2D4_VMS_L2D4PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L2D4_VMS_L2D4PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L2D4_VMS_L2D4PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L2D4_VMS_L2D4PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L2D4_VMS_L2D4PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L2D4_VMS_L2D4PHI2Z2n6),
.vmstuboutPHI3Z2n1(VMR_L2D4_VMS_L2D4PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L2D4_VMS_L2D4PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L2D4_VMS_L2D4PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L2D4_VMS_L2D4PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L2D4_VMS_L2D4PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L2D4_VMS_L2D4PHI3Z2n6),
.vmstuboutPHI4Z2n1(VMR_L2D4_VMS_L2D4PHI4Z2n1),
.vmstuboutPHI4Z2n2(VMR_L2D4_VMS_L2D4PHI4Z2n2),
.vmstuboutPHI4Z2n3(VMR_L2D4_VMS_L2D4PHI4Z2n3),
.vmstuboutPHI4Z2n4(VMR_L2D4_VMS_L2D4PHI4Z2n4),
.allstuboutn1(VMR_L2D4_AS_L2D4n1),
.allstuboutn2(VMR_L2D4_AS_L2D4n2),
.allstuboutn3(VMR_L2D4_AS_L2D4n3),
.allstuboutn4(VMR_L2D4_AS_L2D4n4),
.vmstuboutPHI1Z1n1_wr_en(VMR_L2D4_VMS_L2D4PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L2D4_VMS_L2D4PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L2D4_VMS_L2D4PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L2D4_VMS_L2D4PHI1Z1n4_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L2D4_VMS_L2D4PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L2D4_VMS_L2D4PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L2D4_VMS_L2D4PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L2D4_VMS_L2D4PHI2Z1n4_wr_en),
.vmstuboutPHI2Z1n5_wr_en(VMR_L2D4_VMS_L2D4PHI2Z1n5_wr_en),
.vmstuboutPHI2Z1n6_wr_en(VMR_L2D4_VMS_L2D4PHI2Z1n6_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L2D4_VMS_L2D4PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L2D4_VMS_L2D4PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L2D4_VMS_L2D4PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L2D4_VMS_L2D4PHI3Z1n4_wr_en),
.vmstuboutPHI3Z1n5_wr_en(VMR_L2D4_VMS_L2D4PHI3Z1n5_wr_en),
.vmstuboutPHI3Z1n6_wr_en(VMR_L2D4_VMS_L2D4PHI3Z1n6_wr_en),
.vmstuboutPHI4Z1n1_wr_en(VMR_L2D4_VMS_L2D4PHI4Z1n1_wr_en),
.vmstuboutPHI4Z1n2_wr_en(VMR_L2D4_VMS_L2D4PHI4Z1n2_wr_en),
.vmstuboutPHI4Z1n3_wr_en(VMR_L2D4_VMS_L2D4PHI4Z1n3_wr_en),
.vmstuboutPHI4Z1n4_wr_en(VMR_L2D4_VMS_L2D4PHI4Z1n4_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L2D4_VMS_L2D4PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L2D4_VMS_L2D4PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L2D4_VMS_L2D4PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L2D4_VMS_L2D4PHI1Z2n4_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L2D4_VMS_L2D4PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L2D4_VMS_L2D4PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L2D4_VMS_L2D4PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L2D4_VMS_L2D4PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L2D4_VMS_L2D4PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L2D4_VMS_L2D4PHI2Z2n6_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L2D4_VMS_L2D4PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L2D4_VMS_L2D4PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L2D4_VMS_L2D4PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L2D4_VMS_L2D4PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L2D4_VMS_L2D4PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L2D4_VMS_L2D4PHI3Z2n6_wr_en),
.vmstuboutPHI4Z2n1_wr_en(VMR_L2D4_VMS_L2D4PHI4Z2n1_wr_en),
.vmstuboutPHI4Z2n2_wr_en(VMR_L2D4_VMS_L2D4PHI4Z2n2_wr_en),
.vmstuboutPHI4Z2n3_wr_en(VMR_L2D4_VMS_L2D4PHI4Z2n3_wr_en),
.vmstuboutPHI4Z2n4_wr_en(VMR_L2D4_VMS_L2D4PHI4Z2n4_wr_en),
.valid_data1(VMR_L2D4_AS_L2D4n1_wr_en),
.valid_data2(VMR_L2D4_AS_L2D4n2_wr_en),
.valid_data3(VMR_L2D4_AS_L2D4n3_wr_en),
.valid_data4(VMR_L2D4_AS_L2D4n4_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b0,1'b0) VMR_L4D3(
.number_in1(SL1_L4D3_VMR_L4D3_number),
.read_add1(SL1_L4D3_VMR_L4D3_read_add),
.stubinLink1(SL1_L4D3_VMR_L4D3),
.number_in2(SL2_L4D3_VMR_L4D3_number),
.read_add2(SL2_L4D3_VMR_L4D3_read_add),
.stubinLink2(SL2_L4D3_VMR_L4D3),
.number_in3(SL3_L4D3_VMR_L4D3_number),
.read_add3(SL3_L4D3_VMR_L4D3_read_add),
.stubinLink3(SL3_L4D3_VMR_L4D3),
.vmstuboutPHI1Z1n1(VMR_L4D3_VMS_L4D3PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L4D3_VMS_L4D3PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L4D3_VMS_L4D3PHI1Z1n3),
.vmstuboutPHI2Z1n1(VMR_L4D3_VMS_L4D3PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L4D3_VMS_L4D3PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L4D3_VMS_L4D3PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L4D3_VMS_L4D3PHI2Z1n4),
.vmstuboutPHI3Z1n1(VMR_L4D3_VMS_L4D3PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L4D3_VMS_L4D3PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L4D3_VMS_L4D3PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L4D3_VMS_L4D3PHI3Z1n4),
.vmstuboutPHI4Z1n1(VMR_L4D3_VMS_L4D3PHI4Z1n1),
.vmstuboutPHI4Z1n2(VMR_L4D3_VMS_L4D3PHI4Z1n2),
.vmstuboutPHI4Z1n3(VMR_L4D3_VMS_L4D3PHI4Z1n3),
.vmstuboutPHI1Z2n1(VMR_L4D3_VMS_L4D3PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L4D3_VMS_L4D3PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L4D3_VMS_L4D3PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L4D3_VMS_L4D3PHI1Z2n4),
.vmstuboutPHI2Z2n1(VMR_L4D3_VMS_L4D3PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L4D3_VMS_L4D3PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L4D3_VMS_L4D3PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L4D3_VMS_L4D3PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L4D3_VMS_L4D3PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L4D3_VMS_L4D3PHI2Z2n6),
.vmstuboutPHI3Z2n1(VMR_L4D3_VMS_L4D3PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L4D3_VMS_L4D3PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L4D3_VMS_L4D3PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L4D3_VMS_L4D3PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L4D3_VMS_L4D3PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L4D3_VMS_L4D3PHI3Z2n6),
.vmstuboutPHI4Z2n1(VMR_L4D3_VMS_L4D3PHI4Z2n1),
.vmstuboutPHI4Z2n2(VMR_L4D3_VMS_L4D3PHI4Z2n2),
.vmstuboutPHI4Z2n3(VMR_L4D3_VMS_L4D3PHI4Z2n3),
.vmstuboutPHI4Z2n4(VMR_L4D3_VMS_L4D3PHI4Z2n4),
.allstuboutn1(VMR_L4D3_AS_L4D3n1),
.allstuboutn2(VMR_L4D3_AS_L4D3n2),
.allstuboutn3(VMR_L4D3_AS_L4D3n3),
.vmstuboutPHI1Z1n1_wr_en(VMR_L4D3_VMS_L4D3PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L4D3_VMS_L4D3PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L4D3_VMS_L4D3PHI1Z1n3_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L4D3_VMS_L4D3PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L4D3_VMS_L4D3PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L4D3_VMS_L4D3PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L4D3_VMS_L4D3PHI2Z1n4_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L4D3_VMS_L4D3PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L4D3_VMS_L4D3PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L4D3_VMS_L4D3PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L4D3_VMS_L4D3PHI3Z1n4_wr_en),
.vmstuboutPHI4Z1n1_wr_en(VMR_L4D3_VMS_L4D3PHI4Z1n1_wr_en),
.vmstuboutPHI4Z1n2_wr_en(VMR_L4D3_VMS_L4D3PHI4Z1n2_wr_en),
.vmstuboutPHI4Z1n3_wr_en(VMR_L4D3_VMS_L4D3PHI4Z1n3_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L4D3_VMS_L4D3PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L4D3_VMS_L4D3PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L4D3_VMS_L4D3PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L4D3_VMS_L4D3PHI1Z2n4_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L4D3_VMS_L4D3PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L4D3_VMS_L4D3PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L4D3_VMS_L4D3PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L4D3_VMS_L4D3PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L4D3_VMS_L4D3PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L4D3_VMS_L4D3PHI2Z2n6_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L4D3_VMS_L4D3PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L4D3_VMS_L4D3PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L4D3_VMS_L4D3PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L4D3_VMS_L4D3PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L4D3_VMS_L4D3PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L4D3_VMS_L4D3PHI3Z2n6_wr_en),
.vmstuboutPHI4Z2n1_wr_en(VMR_L4D3_VMS_L4D3PHI4Z2n1_wr_en),
.vmstuboutPHI4Z2n2_wr_en(VMR_L4D3_VMS_L4D3PHI4Z2n2_wr_en),
.vmstuboutPHI4Z2n3_wr_en(VMR_L4D3_VMS_L4D3PHI4Z2n3_wr_en),
.vmstuboutPHI4Z2n4_wr_en(VMR_L4D3_VMS_L4D3PHI4Z2n4_wr_en),
.valid_data1(VMR_L4D3_AS_L4D3n1_wr_en),
.valid_data2(VMR_L4D3_AS_L4D3n2_wr_en),
.valid_data3(VMR_L4D3_AS_L4D3n3_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b0,1'b0) VMR_L4D4(
.number_in1(SL1_L4D4_VMR_L4D4_number),
.read_add1(SL1_L4D4_VMR_L4D4_read_add),
.stubinLink1(SL1_L4D4_VMR_L4D4),
.number_in2(SL2_L4D4_VMR_L4D4_number),
.read_add2(SL2_L4D4_VMR_L4D4_read_add),
.stubinLink2(SL2_L4D4_VMR_L4D4),
.number_in3(SL3_L4D4_VMR_L4D4_number),
.read_add3(SL3_L4D4_VMR_L4D4_read_add),
.stubinLink3(SL3_L4D4_VMR_L4D4),
.vmstuboutPHI1Z1n1(VMR_L4D4_VMS_L4D4PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L4D4_VMS_L4D4PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L4D4_VMS_L4D4PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L4D4_VMS_L4D4PHI1Z1n4),
.vmstuboutPHI2Z1n1(VMR_L4D4_VMS_L4D4PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L4D4_VMS_L4D4PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L4D4_VMS_L4D4PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L4D4_VMS_L4D4PHI2Z1n4),
.vmstuboutPHI2Z1n5(VMR_L4D4_VMS_L4D4PHI2Z1n5),
.vmstuboutPHI2Z1n6(VMR_L4D4_VMS_L4D4PHI2Z1n6),
.vmstuboutPHI3Z1n1(VMR_L4D4_VMS_L4D4PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L4D4_VMS_L4D4PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L4D4_VMS_L4D4PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L4D4_VMS_L4D4PHI3Z1n4),
.vmstuboutPHI3Z1n5(VMR_L4D4_VMS_L4D4PHI3Z1n5),
.vmstuboutPHI3Z1n6(VMR_L4D4_VMS_L4D4PHI3Z1n6),
.vmstuboutPHI4Z1n1(VMR_L4D4_VMS_L4D4PHI4Z1n1),
.vmstuboutPHI4Z1n2(VMR_L4D4_VMS_L4D4PHI4Z1n2),
.vmstuboutPHI4Z1n3(VMR_L4D4_VMS_L4D4PHI4Z1n3),
.vmstuboutPHI4Z1n4(VMR_L4D4_VMS_L4D4PHI4Z1n4),
.vmstuboutPHI1Z2n1(VMR_L4D4_VMS_L4D4PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L4D4_VMS_L4D4PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L4D4_VMS_L4D4PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L4D4_VMS_L4D4PHI1Z2n4),
.vmstuboutPHI2Z2n1(VMR_L4D4_VMS_L4D4PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L4D4_VMS_L4D4PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L4D4_VMS_L4D4PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L4D4_VMS_L4D4PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L4D4_VMS_L4D4PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L4D4_VMS_L4D4PHI2Z2n6),
.vmstuboutPHI3Z2n1(VMR_L4D4_VMS_L4D4PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L4D4_VMS_L4D4PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L4D4_VMS_L4D4PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L4D4_VMS_L4D4PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L4D4_VMS_L4D4PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L4D4_VMS_L4D4PHI3Z2n6),
.vmstuboutPHI4Z2n1(VMR_L4D4_VMS_L4D4PHI4Z2n1),
.vmstuboutPHI4Z2n2(VMR_L4D4_VMS_L4D4PHI4Z2n2),
.vmstuboutPHI4Z2n3(VMR_L4D4_VMS_L4D4PHI4Z2n3),
.vmstuboutPHI4Z2n4(VMR_L4D4_VMS_L4D4PHI4Z2n4),
.allstuboutn1(VMR_L4D4_AS_L4D4n1),
.allstuboutn2(VMR_L4D4_AS_L4D4n2),
.allstuboutn3(VMR_L4D4_AS_L4D4n3),
.allstuboutn4(VMR_L4D4_AS_L4D4n4),
.vmstuboutPHI1Z1n1_wr_en(VMR_L4D4_VMS_L4D4PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L4D4_VMS_L4D4PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L4D4_VMS_L4D4PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L4D4_VMS_L4D4PHI1Z1n4_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L4D4_VMS_L4D4PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L4D4_VMS_L4D4PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L4D4_VMS_L4D4PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L4D4_VMS_L4D4PHI2Z1n4_wr_en),
.vmstuboutPHI2Z1n5_wr_en(VMR_L4D4_VMS_L4D4PHI2Z1n5_wr_en),
.vmstuboutPHI2Z1n6_wr_en(VMR_L4D4_VMS_L4D4PHI2Z1n6_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L4D4_VMS_L4D4PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L4D4_VMS_L4D4PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L4D4_VMS_L4D4PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L4D4_VMS_L4D4PHI3Z1n4_wr_en),
.vmstuboutPHI3Z1n5_wr_en(VMR_L4D4_VMS_L4D4PHI3Z1n5_wr_en),
.vmstuboutPHI3Z1n6_wr_en(VMR_L4D4_VMS_L4D4PHI3Z1n6_wr_en),
.vmstuboutPHI4Z1n1_wr_en(VMR_L4D4_VMS_L4D4PHI4Z1n1_wr_en),
.vmstuboutPHI4Z1n2_wr_en(VMR_L4D4_VMS_L4D4PHI4Z1n2_wr_en),
.vmstuboutPHI4Z1n3_wr_en(VMR_L4D4_VMS_L4D4PHI4Z1n3_wr_en),
.vmstuboutPHI4Z1n4_wr_en(VMR_L4D4_VMS_L4D4PHI4Z1n4_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L4D4_VMS_L4D4PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L4D4_VMS_L4D4PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L4D4_VMS_L4D4PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L4D4_VMS_L4D4PHI1Z2n4_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L4D4_VMS_L4D4PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L4D4_VMS_L4D4PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L4D4_VMS_L4D4PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L4D4_VMS_L4D4PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L4D4_VMS_L4D4PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L4D4_VMS_L4D4PHI2Z2n6_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L4D4_VMS_L4D4PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L4D4_VMS_L4D4PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L4D4_VMS_L4D4PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L4D4_VMS_L4D4PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L4D4_VMS_L4D4PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L4D4_VMS_L4D4PHI3Z2n6_wr_en),
.vmstuboutPHI4Z2n1_wr_en(VMR_L4D4_VMS_L4D4PHI4Z2n1_wr_en),
.vmstuboutPHI4Z2n2_wr_en(VMR_L4D4_VMS_L4D4PHI4Z2n2_wr_en),
.vmstuboutPHI4Z2n3_wr_en(VMR_L4D4_VMS_L4D4PHI4Z2n3_wr_en),
.vmstuboutPHI4Z2n4_wr_en(VMR_L4D4_VMS_L4D4PHI4Z2n4_wr_en),
.valid_data1(VMR_L4D4_AS_L4D4n1_wr_en),
.valid_data2(VMR_L4D4_AS_L4D4n2_wr_en),
.valid_data3(VMR_L4D4_AS_L4D4n3_wr_en),
.valid_data4(VMR_L4D4_AS_L4D4n4_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b0,1'b0) VMR_L6D3(
.number_in1(SL1_L6D3_VMR_L6D3_number),
.read_add1(SL1_L6D3_VMR_L6D3_read_add),
.stubinLink1(SL1_L6D3_VMR_L6D3),
.number_in2(SL2_L6D3_VMR_L6D3_number),
.read_add2(SL2_L6D3_VMR_L6D3_read_add),
.stubinLink2(SL2_L6D3_VMR_L6D3),
.number_in3(SL3_L6D3_VMR_L6D3_number),
.read_add3(SL3_L6D3_VMR_L6D3_read_add),
.stubinLink3(SL3_L6D3_VMR_L6D3),
.vmstuboutPHI1Z1n1(VMR_L6D3_VMS_L6D3PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L6D3_VMS_L6D3PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L6D3_VMS_L6D3PHI1Z1n3),
.vmstuboutPHI2Z1n1(VMR_L6D3_VMS_L6D3PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L6D3_VMS_L6D3PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L6D3_VMS_L6D3PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L6D3_VMS_L6D3PHI2Z1n4),
.vmstuboutPHI3Z1n1(VMR_L6D3_VMS_L6D3PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L6D3_VMS_L6D3PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L6D3_VMS_L6D3PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L6D3_VMS_L6D3PHI3Z1n4),
.vmstuboutPHI4Z1n1(VMR_L6D3_VMS_L6D3PHI4Z1n1),
.vmstuboutPHI4Z1n2(VMR_L6D3_VMS_L6D3PHI4Z1n2),
.vmstuboutPHI4Z1n3(VMR_L6D3_VMS_L6D3PHI4Z1n3),
.vmstuboutPHI1Z2n1(VMR_L6D3_VMS_L6D3PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L6D3_VMS_L6D3PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L6D3_VMS_L6D3PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L6D3_VMS_L6D3PHI1Z2n4),
.vmstuboutPHI2Z2n1(VMR_L6D3_VMS_L6D3PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L6D3_VMS_L6D3PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L6D3_VMS_L6D3PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L6D3_VMS_L6D3PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L6D3_VMS_L6D3PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L6D3_VMS_L6D3PHI2Z2n6),
.vmstuboutPHI3Z2n1(VMR_L6D3_VMS_L6D3PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L6D3_VMS_L6D3PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L6D3_VMS_L6D3PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L6D3_VMS_L6D3PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L6D3_VMS_L6D3PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L6D3_VMS_L6D3PHI3Z2n6),
.vmstuboutPHI4Z2n1(VMR_L6D3_VMS_L6D3PHI4Z2n1),
.vmstuboutPHI4Z2n2(VMR_L6D3_VMS_L6D3PHI4Z2n2),
.vmstuboutPHI4Z2n3(VMR_L6D3_VMS_L6D3PHI4Z2n3),
.vmstuboutPHI4Z2n4(VMR_L6D3_VMS_L6D3PHI4Z2n4),
.allstuboutn1(VMR_L6D3_AS_L6D3n1),
.allstuboutn2(VMR_L6D3_AS_L6D3n2),
.allstuboutn3(VMR_L6D3_AS_L6D3n3),
.vmstuboutPHI1Z1n1_wr_en(VMR_L6D3_VMS_L6D3PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L6D3_VMS_L6D3PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L6D3_VMS_L6D3PHI1Z1n3_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L6D3_VMS_L6D3PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L6D3_VMS_L6D3PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L6D3_VMS_L6D3PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L6D3_VMS_L6D3PHI2Z1n4_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L6D3_VMS_L6D3PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L6D3_VMS_L6D3PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L6D3_VMS_L6D3PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L6D3_VMS_L6D3PHI3Z1n4_wr_en),
.vmstuboutPHI4Z1n1_wr_en(VMR_L6D3_VMS_L6D3PHI4Z1n1_wr_en),
.vmstuboutPHI4Z1n2_wr_en(VMR_L6D3_VMS_L6D3PHI4Z1n2_wr_en),
.vmstuboutPHI4Z1n3_wr_en(VMR_L6D3_VMS_L6D3PHI4Z1n3_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L6D3_VMS_L6D3PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L6D3_VMS_L6D3PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L6D3_VMS_L6D3PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L6D3_VMS_L6D3PHI1Z2n4_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L6D3_VMS_L6D3PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L6D3_VMS_L6D3PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L6D3_VMS_L6D3PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L6D3_VMS_L6D3PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L6D3_VMS_L6D3PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L6D3_VMS_L6D3PHI2Z2n6_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L6D3_VMS_L6D3PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L6D3_VMS_L6D3PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L6D3_VMS_L6D3PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L6D3_VMS_L6D3PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L6D3_VMS_L6D3PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L6D3_VMS_L6D3PHI3Z2n6_wr_en),
.vmstuboutPHI4Z2n1_wr_en(VMR_L6D3_VMS_L6D3PHI4Z2n1_wr_en),
.vmstuboutPHI4Z2n2_wr_en(VMR_L6D3_VMS_L6D3PHI4Z2n2_wr_en),
.vmstuboutPHI4Z2n3_wr_en(VMR_L6D3_VMS_L6D3PHI4Z2n3_wr_en),
.vmstuboutPHI4Z2n4_wr_en(VMR_L6D3_VMS_L6D3PHI4Z2n4_wr_en),
.valid_data1(VMR_L6D3_AS_L6D3n1_wr_en),
.valid_data2(VMR_L6D3_AS_L6D3n2_wr_en),
.valid_data3(VMR_L6D3_AS_L6D3n3_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


VMRouter #(1'b0,1'b0) VMR_L6D4(
.number_in1(SL1_L6D4_VMR_L6D4_number),
.read_add1(SL1_L6D4_VMR_L6D4_read_add),
.stubinLink1(SL1_L6D4_VMR_L6D4),
.number_in2(SL2_L6D4_VMR_L6D4_number),
.read_add2(SL2_L6D4_VMR_L6D4_read_add),
.stubinLink2(SL2_L6D4_VMR_L6D4),
.number_in3(SL3_L6D4_VMR_L6D4_number),
.read_add3(SL3_L6D4_VMR_L6D4_read_add),
.stubinLink3(SL3_L6D4_VMR_L6D4),
.vmstuboutPHI1Z1n1(VMR_L6D4_VMS_L6D4PHI1Z1n1),
.vmstuboutPHI1Z1n2(VMR_L6D4_VMS_L6D4PHI1Z1n2),
.vmstuboutPHI1Z1n3(VMR_L6D4_VMS_L6D4PHI1Z1n3),
.vmstuboutPHI1Z1n4(VMR_L6D4_VMS_L6D4PHI1Z1n4),
.vmstuboutPHI2Z1n1(VMR_L6D4_VMS_L6D4PHI2Z1n1),
.vmstuboutPHI2Z1n2(VMR_L6D4_VMS_L6D4PHI2Z1n2),
.vmstuboutPHI2Z1n3(VMR_L6D4_VMS_L6D4PHI2Z1n3),
.vmstuboutPHI2Z1n4(VMR_L6D4_VMS_L6D4PHI2Z1n4),
.vmstuboutPHI2Z1n5(VMR_L6D4_VMS_L6D4PHI2Z1n5),
.vmstuboutPHI2Z1n6(VMR_L6D4_VMS_L6D4PHI2Z1n6),
.vmstuboutPHI3Z1n1(VMR_L6D4_VMS_L6D4PHI3Z1n1),
.vmstuboutPHI3Z1n2(VMR_L6D4_VMS_L6D4PHI3Z1n2),
.vmstuboutPHI3Z1n3(VMR_L6D4_VMS_L6D4PHI3Z1n3),
.vmstuboutPHI3Z1n4(VMR_L6D4_VMS_L6D4PHI3Z1n4),
.vmstuboutPHI3Z1n5(VMR_L6D4_VMS_L6D4PHI3Z1n5),
.vmstuboutPHI3Z1n6(VMR_L6D4_VMS_L6D4PHI3Z1n6),
.vmstuboutPHI4Z1n1(VMR_L6D4_VMS_L6D4PHI4Z1n1),
.vmstuboutPHI4Z1n2(VMR_L6D4_VMS_L6D4PHI4Z1n2),
.vmstuboutPHI4Z1n3(VMR_L6D4_VMS_L6D4PHI4Z1n3),
.vmstuboutPHI4Z1n4(VMR_L6D4_VMS_L6D4PHI4Z1n4),
.vmstuboutPHI1Z2n1(VMR_L6D4_VMS_L6D4PHI1Z2n1),
.vmstuboutPHI1Z2n2(VMR_L6D4_VMS_L6D4PHI1Z2n2),
.vmstuboutPHI1Z2n3(VMR_L6D4_VMS_L6D4PHI1Z2n3),
.vmstuboutPHI1Z2n4(VMR_L6D4_VMS_L6D4PHI1Z2n4),
.vmstuboutPHI2Z2n1(VMR_L6D4_VMS_L6D4PHI2Z2n1),
.vmstuboutPHI2Z2n2(VMR_L6D4_VMS_L6D4PHI2Z2n2),
.vmstuboutPHI2Z2n3(VMR_L6D4_VMS_L6D4PHI2Z2n3),
.vmstuboutPHI2Z2n4(VMR_L6D4_VMS_L6D4PHI2Z2n4),
.vmstuboutPHI2Z2n5(VMR_L6D4_VMS_L6D4PHI2Z2n5),
.vmstuboutPHI2Z2n6(VMR_L6D4_VMS_L6D4PHI2Z2n6),
.vmstuboutPHI3Z2n1(VMR_L6D4_VMS_L6D4PHI3Z2n1),
.vmstuboutPHI3Z2n2(VMR_L6D4_VMS_L6D4PHI3Z2n2),
.vmstuboutPHI3Z2n3(VMR_L6D4_VMS_L6D4PHI3Z2n3),
.vmstuboutPHI3Z2n4(VMR_L6D4_VMS_L6D4PHI3Z2n4),
.vmstuboutPHI3Z2n5(VMR_L6D4_VMS_L6D4PHI3Z2n5),
.vmstuboutPHI3Z2n6(VMR_L6D4_VMS_L6D4PHI3Z2n6),
.vmstuboutPHI4Z2n1(VMR_L6D4_VMS_L6D4PHI4Z2n1),
.vmstuboutPHI4Z2n2(VMR_L6D4_VMS_L6D4PHI4Z2n2),
.vmstuboutPHI4Z2n3(VMR_L6D4_VMS_L6D4PHI4Z2n3),
.vmstuboutPHI4Z2n4(VMR_L6D4_VMS_L6D4PHI4Z2n4),
.allstuboutn1(VMR_L6D4_AS_L6D4n1),
.allstuboutn2(VMR_L6D4_AS_L6D4n2),
.allstuboutn3(VMR_L6D4_AS_L6D4n3),
.allstuboutn4(VMR_L6D4_AS_L6D4n4),
.vmstuboutPHI1Z1n1_wr_en(VMR_L6D4_VMS_L6D4PHI1Z1n1_wr_en),
.vmstuboutPHI1Z1n2_wr_en(VMR_L6D4_VMS_L6D4PHI1Z1n2_wr_en),
.vmstuboutPHI1Z1n3_wr_en(VMR_L6D4_VMS_L6D4PHI1Z1n3_wr_en),
.vmstuboutPHI1Z1n4_wr_en(VMR_L6D4_VMS_L6D4PHI1Z1n4_wr_en),
.vmstuboutPHI2Z1n1_wr_en(VMR_L6D4_VMS_L6D4PHI2Z1n1_wr_en),
.vmstuboutPHI2Z1n2_wr_en(VMR_L6D4_VMS_L6D4PHI2Z1n2_wr_en),
.vmstuboutPHI2Z1n3_wr_en(VMR_L6D4_VMS_L6D4PHI2Z1n3_wr_en),
.vmstuboutPHI2Z1n4_wr_en(VMR_L6D4_VMS_L6D4PHI2Z1n4_wr_en),
.vmstuboutPHI2Z1n5_wr_en(VMR_L6D4_VMS_L6D4PHI2Z1n5_wr_en),
.vmstuboutPHI2Z1n6_wr_en(VMR_L6D4_VMS_L6D4PHI2Z1n6_wr_en),
.vmstuboutPHI3Z1n1_wr_en(VMR_L6D4_VMS_L6D4PHI3Z1n1_wr_en),
.vmstuboutPHI3Z1n2_wr_en(VMR_L6D4_VMS_L6D4PHI3Z1n2_wr_en),
.vmstuboutPHI3Z1n3_wr_en(VMR_L6D4_VMS_L6D4PHI3Z1n3_wr_en),
.vmstuboutPHI3Z1n4_wr_en(VMR_L6D4_VMS_L6D4PHI3Z1n4_wr_en),
.vmstuboutPHI3Z1n5_wr_en(VMR_L6D4_VMS_L6D4PHI3Z1n5_wr_en),
.vmstuboutPHI3Z1n6_wr_en(VMR_L6D4_VMS_L6D4PHI3Z1n6_wr_en),
.vmstuboutPHI4Z1n1_wr_en(VMR_L6D4_VMS_L6D4PHI4Z1n1_wr_en),
.vmstuboutPHI4Z1n2_wr_en(VMR_L6D4_VMS_L6D4PHI4Z1n2_wr_en),
.vmstuboutPHI4Z1n3_wr_en(VMR_L6D4_VMS_L6D4PHI4Z1n3_wr_en),
.vmstuboutPHI4Z1n4_wr_en(VMR_L6D4_VMS_L6D4PHI4Z1n4_wr_en),
.vmstuboutPHI1Z2n1_wr_en(VMR_L6D4_VMS_L6D4PHI1Z2n1_wr_en),
.vmstuboutPHI1Z2n2_wr_en(VMR_L6D4_VMS_L6D4PHI1Z2n2_wr_en),
.vmstuboutPHI1Z2n3_wr_en(VMR_L6D4_VMS_L6D4PHI1Z2n3_wr_en),
.vmstuboutPHI1Z2n4_wr_en(VMR_L6D4_VMS_L6D4PHI1Z2n4_wr_en),
.vmstuboutPHI2Z2n1_wr_en(VMR_L6D4_VMS_L6D4PHI2Z2n1_wr_en),
.vmstuboutPHI2Z2n2_wr_en(VMR_L6D4_VMS_L6D4PHI2Z2n2_wr_en),
.vmstuboutPHI2Z2n3_wr_en(VMR_L6D4_VMS_L6D4PHI2Z2n3_wr_en),
.vmstuboutPHI2Z2n4_wr_en(VMR_L6D4_VMS_L6D4PHI2Z2n4_wr_en),
.vmstuboutPHI2Z2n5_wr_en(VMR_L6D4_VMS_L6D4PHI2Z2n5_wr_en),
.vmstuboutPHI2Z2n6_wr_en(VMR_L6D4_VMS_L6D4PHI2Z2n6_wr_en),
.vmstuboutPHI3Z2n1_wr_en(VMR_L6D4_VMS_L6D4PHI3Z2n1_wr_en),
.vmstuboutPHI3Z2n2_wr_en(VMR_L6D4_VMS_L6D4PHI3Z2n2_wr_en),
.vmstuboutPHI3Z2n3_wr_en(VMR_L6D4_VMS_L6D4PHI3Z2n3_wr_en),
.vmstuboutPHI3Z2n4_wr_en(VMR_L6D4_VMS_L6D4PHI3Z2n4_wr_en),
.vmstuboutPHI3Z2n5_wr_en(VMR_L6D4_VMS_L6D4PHI3Z2n5_wr_en),
.vmstuboutPHI3Z2n6_wr_en(VMR_L6D4_VMS_L6D4PHI3Z2n6_wr_en),
.vmstuboutPHI4Z2n1_wr_en(VMR_L6D4_VMS_L6D4PHI4Z2n1_wr_en),
.vmstuboutPHI4Z2n2_wr_en(VMR_L6D4_VMS_L6D4PHI4Z2n2_wr_en),
.vmstuboutPHI4Z2n3_wr_en(VMR_L6D4_VMS_L6D4PHI4Z2n3_wr_en),
.vmstuboutPHI4Z2n4_wr_en(VMR_L6D4_VMS_L6D4PHI4Z2n4_wr_en),
.valid_data1(VMR_L6D4_AS_L6D4n1_wr_en),
.valid_data2(VMR_L6D4_AS_L6D4n2_wr_en),
.valid_data3(VMR_L6D4_AS_L6D4n3_wr_en),
.valid_data4(VMR_L6D4_AS_L6D4n4_wr_en),
.start(start2_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z1_L2D3PHI1Z1_phi.txt","TETable_TE_L1D3PHI1Z1_L2D3PHI1Z1_z.txt") TE_L1D3PHI1Z1_L2D3PHI1Z1(
.number_in1(VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_number),
.read_add1(VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_read_add),
.innervmstubin(VMS_L1D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1),
.number_in2(VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_number),
.read_add2(VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1_read_add),
.outervmstubin(VMS_L2D3PHI1Z1n1_TE_L1D3PHI1Z1_L2D3PHI1Z1),
.stubpairout(TE_L1D3PHI1Z1_L2D3PHI1Z1_SP_L1D3PHI1Z1_L2D3PHI1Z1),
.valid_data(TE_L1D3PHI1Z1_L2D3PHI1Z1_SP_L1D3PHI1Z1_L2D3PHI1Z1_wr_en),
.start(start3_5),
.done(done3_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z1_L2D3PHI2Z1_phi.txt","TETable_TE_L1D3PHI1Z1_L2D3PHI2Z1_z.txt") TE_L1D3PHI1Z1_L2D3PHI2Z1(
.number_in1(VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1_number),
.read_add1(VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1_read_add),
.innervmstubin(VMS_L1D3PHI1Z1n2_TE_L1D3PHI1Z1_L2D3PHI2Z1),
.number_in2(VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1_number),
.read_add2(VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1_read_add),
.outervmstubin(VMS_L2D3PHI2Z1n1_TE_L1D3PHI1Z1_L2D3PHI2Z1),
.stubpairout(TE_L1D3PHI1Z1_L2D3PHI2Z1_SP_L1D3PHI1Z1_L2D3PHI2Z1),
.valid_data(TE_L1D3PHI1Z1_L2D3PHI2Z1_SP_L1D3PHI1Z1_L2D3PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z1_L2D3PHI2Z1_phi.txt","TETable_TE_L1D3PHI2Z1_L2D3PHI2Z1_z.txt") TE_L1D3PHI2Z1_L2D3PHI2Z1(
.number_in1(VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1_number),
.read_add1(VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1_read_add),
.outervmstubin(VMS_L2D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI2Z1),
.number_in2(VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1_number),
.read_add2(VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1_read_add),
.innervmstubin(VMS_L1D3PHI2Z1n1_TE_L1D3PHI2Z1_L2D3PHI2Z1),
.stubpairout(TE_L1D3PHI2Z1_L2D3PHI2Z1_SP_L1D3PHI2Z1_L2D3PHI2Z1),
.valid_data(TE_L1D3PHI2Z1_L2D3PHI2Z1_SP_L1D3PHI2Z1_L2D3PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z1_L2D3PHI3Z1_phi.txt","TETable_TE_L1D3PHI2Z1_L2D3PHI3Z1_z.txt") TE_L1D3PHI2Z1_L2D3PHI3Z1(
.number_in1(VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1_number),
.read_add1(VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1_read_add),
.innervmstubin(VMS_L1D3PHI2Z1n2_TE_L1D3PHI2Z1_L2D3PHI3Z1),
.number_in2(VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1_number),
.read_add2(VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1_read_add),
.outervmstubin(VMS_L2D3PHI3Z1n1_TE_L1D3PHI2Z1_L2D3PHI3Z1),
.stubpairout(TE_L1D3PHI2Z1_L2D3PHI3Z1_SP_L1D3PHI2Z1_L2D3PHI3Z1),
.valid_data(TE_L1D3PHI2Z1_L2D3PHI3Z1_SP_L1D3PHI2Z1_L2D3PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z1_L2D3PHI3Z1_phi.txt","TETable_TE_L1D3PHI3Z1_L2D3PHI3Z1_z.txt") TE_L1D3PHI3Z1_L2D3PHI3Z1(
.number_in1(VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1_number),
.read_add1(VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1_read_add),
.outervmstubin(VMS_L2D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI3Z1),
.number_in2(VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1_number),
.read_add2(VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1_read_add),
.innervmstubin(VMS_L1D3PHI3Z1n1_TE_L1D3PHI3Z1_L2D3PHI3Z1),
.stubpairout(TE_L1D3PHI3Z1_L2D3PHI3Z1_SP_L1D3PHI3Z1_L2D3PHI3Z1),
.valid_data(TE_L1D3PHI3Z1_L2D3PHI3Z1_SP_L1D3PHI3Z1_L2D3PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z1_L2D3PHI4Z1_phi.txt","TETable_TE_L1D3PHI3Z1_L2D3PHI4Z1_z.txt") TE_L1D3PHI3Z1_L2D3PHI4Z1(
.number_in1(VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1_number),
.read_add1(VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1_read_add),
.innervmstubin(VMS_L1D3PHI3Z1n2_TE_L1D3PHI3Z1_L2D3PHI4Z1),
.number_in2(VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1_number),
.read_add2(VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1_read_add),
.outervmstubin(VMS_L2D3PHI4Z1n1_TE_L1D3PHI3Z1_L2D3PHI4Z1),
.stubpairout(TE_L1D3PHI3Z1_L2D3PHI4Z1_SP_L1D3PHI3Z1_L2D3PHI4Z1),
.valid_data(TE_L1D3PHI3Z1_L2D3PHI4Z1_SP_L1D3PHI3Z1_L2D3PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z1_L2D3PHI1Z2_phi.txt","TETable_TE_L1D3PHI1Z1_L2D3PHI1Z2_z.txt") TE_L1D3PHI1Z1_L2D3PHI1Z2(
.number_in1(VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2_number),
.read_add1(VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2_read_add),
.innervmstubin(VMS_L1D3PHI1Z1n3_TE_L1D3PHI1Z1_L2D3PHI1Z2),
.number_in2(VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2_number),
.read_add2(VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2_read_add),
.outervmstubin(VMS_L2D3PHI1Z2n1_TE_L1D3PHI1Z1_L2D3PHI1Z2),
.stubpairout(TE_L1D3PHI1Z1_L2D3PHI1Z2_SP_L1D3PHI1Z1_L2D3PHI1Z2),
.valid_data(TE_L1D3PHI1Z1_L2D3PHI1Z2_SP_L1D3PHI1Z1_L2D3PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z1_L2D3PHI2Z2_phi.txt","TETable_TE_L1D3PHI1Z1_L2D3PHI2Z2_z.txt") TE_L1D3PHI1Z1_L2D3PHI2Z2(
.number_in1(VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2_number),
.read_add1(VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2_read_add),
.innervmstubin(VMS_L1D3PHI1Z1n4_TE_L1D3PHI1Z1_L2D3PHI2Z2),
.number_in2(VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2_number),
.read_add2(VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2_read_add),
.outervmstubin(VMS_L2D3PHI2Z2n1_TE_L1D3PHI1Z1_L2D3PHI2Z2),
.stubpairout(TE_L1D3PHI1Z1_L2D3PHI2Z2_SP_L1D3PHI1Z1_L2D3PHI2Z2),
.valid_data(TE_L1D3PHI1Z1_L2D3PHI2Z2_SP_L1D3PHI1Z1_L2D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z1_L2D3PHI2Z2_phi.txt","TETable_TE_L1D3PHI2Z1_L2D3PHI2Z2_z.txt") TE_L1D3PHI2Z1_L2D3PHI2Z2(
.number_in1(VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2_number),
.read_add1(VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2_read_add),
.innervmstubin(VMS_L1D3PHI2Z1n3_TE_L1D3PHI2Z1_L2D3PHI2Z2),
.number_in2(VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2_number),
.read_add2(VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2_read_add),
.outervmstubin(VMS_L2D3PHI2Z2n2_TE_L1D3PHI2Z1_L2D3PHI2Z2),
.stubpairout(TE_L1D3PHI2Z1_L2D3PHI2Z2_SP_L1D3PHI2Z1_L2D3PHI2Z2),
.valid_data(TE_L1D3PHI2Z1_L2D3PHI2Z2_SP_L1D3PHI2Z1_L2D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z1_L2D3PHI3Z2_phi.txt","TETable_TE_L1D3PHI2Z1_L2D3PHI3Z2_z.txt") TE_L1D3PHI2Z1_L2D3PHI3Z2(
.number_in1(VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2_number),
.read_add1(VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2_read_add),
.innervmstubin(VMS_L1D3PHI2Z1n4_TE_L1D3PHI2Z1_L2D3PHI3Z2),
.number_in2(VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2_number),
.read_add2(VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2_read_add),
.outervmstubin(VMS_L2D3PHI3Z2n1_TE_L1D3PHI2Z1_L2D3PHI3Z2),
.stubpairout(TE_L1D3PHI2Z1_L2D3PHI3Z2_SP_L1D3PHI2Z1_L2D3PHI3Z2),
.valid_data(TE_L1D3PHI2Z1_L2D3PHI3Z2_SP_L1D3PHI2Z1_L2D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z1_L2D3PHI3Z2_phi.txt","TETable_TE_L1D3PHI3Z1_L2D3PHI3Z2_z.txt") TE_L1D3PHI3Z1_L2D3PHI3Z2(
.number_in1(VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2_number),
.read_add1(VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2_read_add),
.innervmstubin(VMS_L1D3PHI3Z1n3_TE_L1D3PHI3Z1_L2D3PHI3Z2),
.number_in2(VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2_number),
.read_add2(VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2_read_add),
.outervmstubin(VMS_L2D3PHI3Z2n2_TE_L1D3PHI3Z1_L2D3PHI3Z2),
.stubpairout(TE_L1D3PHI3Z1_L2D3PHI3Z2_SP_L1D3PHI3Z1_L2D3PHI3Z2),
.valid_data(TE_L1D3PHI3Z1_L2D3PHI3Z2_SP_L1D3PHI3Z1_L2D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z1_L2D3PHI4Z2_phi.txt","TETable_TE_L1D3PHI3Z1_L2D3PHI4Z2_z.txt") TE_L1D3PHI3Z1_L2D3PHI4Z2(
.number_in1(VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2_number),
.read_add1(VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2_read_add),
.innervmstubin(VMS_L1D3PHI3Z1n4_TE_L1D3PHI3Z1_L2D3PHI4Z2),
.number_in2(VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2_number),
.read_add2(VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2_read_add),
.outervmstubin(VMS_L2D3PHI4Z2n1_TE_L1D3PHI3Z1_L2D3PHI4Z2),
.stubpairout(TE_L1D3PHI3Z1_L2D3PHI4Z2_SP_L1D3PHI3Z1_L2D3PHI4Z2),
.valid_data(TE_L1D3PHI3Z1_L2D3PHI4Z2_SP_L1D3PHI3Z1_L2D3PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z2_L2D3PHI1Z2_phi.txt","TETable_TE_L1D3PHI1Z2_L2D3PHI1Z2_z.txt") TE_L1D3PHI1Z2_L2D3PHI1Z2(
.number_in1(VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2_number),
.read_add1(VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2_read_add),
.outervmstubin(VMS_L2D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI1Z2),
.number_in2(VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2_number),
.read_add2(VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2_read_add),
.innervmstubin(VMS_L1D3PHI1Z2n1_TE_L1D3PHI1Z2_L2D3PHI1Z2),
.stubpairout(TE_L1D3PHI1Z2_L2D3PHI1Z2_SP_L1D3PHI1Z2_L2D3PHI1Z2),
.valid_data(TE_L1D3PHI1Z2_L2D3PHI1Z2_SP_L1D3PHI1Z2_L2D3PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z2_L2D3PHI2Z2_phi.txt","TETable_TE_L1D3PHI1Z2_L2D3PHI2Z2_z.txt") TE_L1D3PHI1Z2_L2D3PHI2Z2(
.number_in1(VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2_number),
.read_add1(VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2_read_add),
.outervmstubin(VMS_L2D3PHI2Z2n3_TE_L1D3PHI1Z2_L2D3PHI2Z2),
.number_in2(VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2_number),
.read_add2(VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2_read_add),
.innervmstubin(VMS_L1D3PHI1Z2n2_TE_L1D3PHI1Z2_L2D3PHI2Z2),
.stubpairout(TE_L1D3PHI1Z2_L2D3PHI2Z2_SP_L1D3PHI1Z2_L2D3PHI2Z2),
.valid_data(TE_L1D3PHI1Z2_L2D3PHI2Z2_SP_L1D3PHI1Z2_L2D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z2_L2D3PHI2Z2_phi.txt","TETable_TE_L1D3PHI2Z2_L2D3PHI2Z2_z.txt") TE_L1D3PHI2Z2_L2D3PHI2Z2(
.number_in1(VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2_number),
.read_add1(VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2_read_add),
.outervmstubin(VMS_L2D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D3PHI2Z2),
.number_in2(VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2_number),
.read_add2(VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2_read_add),
.innervmstubin(VMS_L1D3PHI2Z2n1_TE_L1D3PHI2Z2_L2D3PHI2Z2),
.stubpairout(TE_L1D3PHI2Z2_L2D3PHI2Z2_SP_L1D3PHI2Z2_L2D3PHI2Z2),
.valid_data(TE_L1D3PHI2Z2_L2D3PHI2Z2_SP_L1D3PHI2Z2_L2D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z2_L2D3PHI3Z2_phi.txt","TETable_TE_L1D3PHI2Z2_L2D3PHI3Z2_z.txt") TE_L1D3PHI2Z2_L2D3PHI3Z2(
.number_in1(VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2_number),
.read_add1(VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2_read_add),
.outervmstubin(VMS_L2D3PHI3Z2n3_TE_L1D3PHI2Z2_L2D3PHI3Z2),
.number_in2(VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2_number),
.read_add2(VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2_read_add),
.innervmstubin(VMS_L1D3PHI2Z2n2_TE_L1D3PHI2Z2_L2D3PHI3Z2),
.stubpairout(TE_L1D3PHI2Z2_L2D3PHI3Z2_SP_L1D3PHI2Z2_L2D3PHI3Z2),
.valid_data(TE_L1D3PHI2Z2_L2D3PHI3Z2_SP_L1D3PHI2Z2_L2D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z2_L2D3PHI3Z2_phi.txt","TETable_TE_L1D3PHI3Z2_L2D3PHI3Z2_z.txt") TE_L1D3PHI3Z2_L2D3PHI3Z2(
.number_in1(VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2_number),
.read_add1(VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2_read_add),
.outervmstubin(VMS_L2D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D3PHI3Z2),
.number_in2(VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2_number),
.read_add2(VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2_read_add),
.innervmstubin(VMS_L1D3PHI3Z2n1_TE_L1D3PHI3Z2_L2D3PHI3Z2),
.stubpairout(TE_L1D3PHI3Z2_L2D3PHI3Z2_SP_L1D3PHI3Z2_L2D3PHI3Z2),
.valid_data(TE_L1D3PHI3Z2_L2D3PHI3Z2_SP_L1D3PHI3Z2_L2D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z2_L2D3PHI4Z2_phi.txt","TETable_TE_L1D3PHI3Z2_L2D3PHI4Z2_z.txt") TE_L1D3PHI3Z2_L2D3PHI4Z2(
.number_in1(VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_number),
.read_add1(VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_read_add),
.outervmstubin(VMS_L2D3PHI4Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2),
.number_in2(VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_number),
.read_add2(VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2_read_add),
.innervmstubin(VMS_L1D3PHI3Z2n2_TE_L1D3PHI3Z2_L2D3PHI4Z2),
.stubpairout(TE_L1D3PHI3Z2_L2D3PHI4Z2_SP_L1D3PHI3Z2_L2D3PHI4Z2),
.valid_data(TE_L1D3PHI3Z2_L2D3PHI4Z2_SP_L1D3PHI3Z2_L2D3PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z1_L2D4PHI1Z1_phi.txt","TETable_TE_L1D3PHI1Z1_L2D4PHI1Z1_z.txt") TE_L1D3PHI1Z1_L2D4PHI1Z1(
.number_in1(VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1_number),
.read_add1(VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1_read_add),
.innervmstubin(VMS_L1D3PHI1Z1n5_TE_L1D3PHI1Z1_L2D4PHI1Z1),
.number_in2(VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1_number),
.read_add2(VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1_read_add),
.outervmstubin(VMS_L2D4PHI1Z1n1_TE_L1D3PHI1Z1_L2D4PHI1Z1),
.stubpairout(TE_L1D3PHI1Z1_L2D4PHI1Z1_SP_L1D3PHI1Z1_L2D4PHI1Z1),
.valid_data(TE_L1D3PHI1Z1_L2D4PHI1Z1_SP_L1D3PHI1Z1_L2D4PHI1Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z1_L2D4PHI2Z1_phi.txt","TETable_TE_L1D3PHI1Z1_L2D4PHI2Z1_z.txt") TE_L1D3PHI1Z1_L2D4PHI2Z1(
.number_in1(VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1_number),
.read_add1(VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1_read_add),
.innervmstubin(VMS_L1D3PHI1Z1n6_TE_L1D3PHI1Z1_L2D4PHI2Z1),
.number_in2(VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1_number),
.read_add2(VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1_read_add),
.outervmstubin(VMS_L2D4PHI2Z1n1_TE_L1D3PHI1Z1_L2D4PHI2Z1),
.stubpairout(TE_L1D3PHI1Z1_L2D4PHI2Z1_SP_L1D3PHI1Z1_L2D4PHI2Z1),
.valid_data(TE_L1D3PHI1Z1_L2D4PHI2Z1_SP_L1D3PHI1Z1_L2D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z1_L2D4PHI2Z1_phi.txt","TETable_TE_L1D3PHI2Z1_L2D4PHI2Z1_z.txt") TE_L1D3PHI2Z1_L2D4PHI2Z1(
.number_in1(VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1_number),
.read_add1(VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1_read_add),
.innervmstubin(VMS_L1D3PHI2Z1n5_TE_L1D3PHI2Z1_L2D4PHI2Z1),
.number_in2(VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1_number),
.read_add2(VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1_read_add),
.outervmstubin(VMS_L2D4PHI2Z1n2_TE_L1D3PHI2Z1_L2D4PHI2Z1),
.stubpairout(TE_L1D3PHI2Z1_L2D4PHI2Z1_SP_L1D3PHI2Z1_L2D4PHI2Z1),
.valid_data(TE_L1D3PHI2Z1_L2D4PHI2Z1_SP_L1D3PHI2Z1_L2D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z1_L2D4PHI3Z1_phi.txt","TETable_TE_L1D3PHI2Z1_L2D4PHI3Z1_z.txt") TE_L1D3PHI2Z1_L2D4PHI3Z1(
.number_in1(VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1_number),
.read_add1(VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1_read_add),
.innervmstubin(VMS_L1D3PHI2Z1n6_TE_L1D3PHI2Z1_L2D4PHI3Z1),
.number_in2(VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1_number),
.read_add2(VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1_read_add),
.outervmstubin(VMS_L2D4PHI3Z1n1_TE_L1D3PHI2Z1_L2D4PHI3Z1),
.stubpairout(TE_L1D3PHI2Z1_L2D4PHI3Z1_SP_L1D3PHI2Z1_L2D4PHI3Z1),
.valid_data(TE_L1D3PHI2Z1_L2D4PHI3Z1_SP_L1D3PHI2Z1_L2D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z1_L2D4PHI3Z1_phi.txt","TETable_TE_L1D3PHI3Z1_L2D4PHI3Z1_z.txt") TE_L1D3PHI3Z1_L2D4PHI3Z1(
.number_in1(VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1_number),
.read_add1(VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1_read_add),
.innervmstubin(VMS_L1D3PHI3Z1n5_TE_L1D3PHI3Z1_L2D4PHI3Z1),
.number_in2(VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1_number),
.read_add2(VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1_read_add),
.outervmstubin(VMS_L2D4PHI3Z1n2_TE_L1D3PHI3Z1_L2D4PHI3Z1),
.stubpairout(TE_L1D3PHI3Z1_L2D4PHI3Z1_SP_L1D3PHI3Z1_L2D4PHI3Z1),
.valid_data(TE_L1D3PHI3Z1_L2D4PHI3Z1_SP_L1D3PHI3Z1_L2D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z1_L2D4PHI4Z1_phi.txt","TETable_TE_L1D3PHI3Z1_L2D4PHI4Z1_z.txt") TE_L1D3PHI3Z1_L2D4PHI4Z1(
.number_in1(VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1_number),
.read_add1(VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1_read_add),
.innervmstubin(VMS_L1D3PHI3Z1n6_TE_L1D3PHI3Z1_L2D4PHI4Z1),
.number_in2(VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1_number),
.read_add2(VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1_read_add),
.outervmstubin(VMS_L2D4PHI4Z1n1_TE_L1D3PHI3Z1_L2D4PHI4Z1),
.stubpairout(TE_L1D3PHI3Z1_L2D4PHI4Z1_SP_L1D3PHI3Z1_L2D4PHI4Z1),
.valid_data(TE_L1D3PHI3Z1_L2D4PHI4Z1_SP_L1D3PHI3Z1_L2D4PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z2_L2D4PHI1Z1_phi.txt","TETable_TE_L1D3PHI1Z2_L2D4PHI1Z1_z.txt") TE_L1D3PHI1Z2_L2D4PHI1Z1(
.number_in1(VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1_number),
.read_add1(VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1_read_add),
.innervmstubin(VMS_L1D3PHI1Z2n3_TE_L1D3PHI1Z2_L2D4PHI1Z1),
.number_in2(VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1_number),
.read_add2(VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1_read_add),
.outervmstubin(VMS_L2D4PHI1Z1n2_TE_L1D3PHI1Z2_L2D4PHI1Z1),
.stubpairout(TE_L1D3PHI1Z2_L2D4PHI1Z1_SP_L1D3PHI1Z2_L2D4PHI1Z1),
.valid_data(TE_L1D3PHI1Z2_L2D4PHI1Z1_SP_L1D3PHI1Z2_L2D4PHI1Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z2_L2D4PHI2Z1_phi.txt","TETable_TE_L1D3PHI1Z2_L2D4PHI2Z1_z.txt") TE_L1D3PHI1Z2_L2D4PHI2Z1(
.number_in1(VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1_number),
.read_add1(VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1_read_add),
.innervmstubin(VMS_L1D3PHI1Z2n4_TE_L1D3PHI1Z2_L2D4PHI2Z1),
.number_in2(VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1_number),
.read_add2(VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1_read_add),
.outervmstubin(VMS_L2D4PHI2Z1n3_TE_L1D3PHI1Z2_L2D4PHI2Z1),
.stubpairout(TE_L1D3PHI1Z2_L2D4PHI2Z1_SP_L1D3PHI1Z2_L2D4PHI2Z1),
.valid_data(TE_L1D3PHI1Z2_L2D4PHI2Z1_SP_L1D3PHI1Z2_L2D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z2_L2D4PHI2Z1_phi.txt","TETable_TE_L1D3PHI2Z2_L2D4PHI2Z1_z.txt") TE_L1D3PHI2Z2_L2D4PHI2Z1(
.number_in1(VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1_number),
.read_add1(VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1_read_add),
.innervmstubin(VMS_L1D3PHI2Z2n3_TE_L1D3PHI2Z2_L2D4PHI2Z1),
.number_in2(VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1_number),
.read_add2(VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1_read_add),
.outervmstubin(VMS_L2D4PHI2Z1n4_TE_L1D3PHI2Z2_L2D4PHI2Z1),
.stubpairout(TE_L1D3PHI2Z2_L2D4PHI2Z1_SP_L1D3PHI2Z2_L2D4PHI2Z1),
.valid_data(TE_L1D3PHI2Z2_L2D4PHI2Z1_SP_L1D3PHI2Z2_L2D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z2_L2D4PHI3Z1_phi.txt","TETable_TE_L1D3PHI2Z2_L2D4PHI3Z1_z.txt") TE_L1D3PHI2Z2_L2D4PHI3Z1(
.number_in1(VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1_number),
.read_add1(VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1_read_add),
.innervmstubin(VMS_L1D3PHI2Z2n4_TE_L1D3PHI2Z2_L2D4PHI3Z1),
.number_in2(VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1_number),
.read_add2(VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1_read_add),
.outervmstubin(VMS_L2D4PHI3Z1n3_TE_L1D3PHI2Z2_L2D4PHI3Z1),
.stubpairout(TE_L1D3PHI2Z2_L2D4PHI3Z1_SP_L1D3PHI2Z2_L2D4PHI3Z1),
.valid_data(TE_L1D3PHI2Z2_L2D4PHI3Z1_SP_L1D3PHI2Z2_L2D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z2_L2D4PHI3Z1_phi.txt","TETable_TE_L1D3PHI3Z2_L2D4PHI3Z1_z.txt") TE_L1D3PHI3Z2_L2D4PHI3Z1(
.number_in1(VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1_number),
.read_add1(VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1_read_add),
.innervmstubin(VMS_L1D3PHI3Z2n3_TE_L1D3PHI3Z2_L2D4PHI3Z1),
.number_in2(VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1_number),
.read_add2(VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1_read_add),
.outervmstubin(VMS_L2D4PHI3Z1n4_TE_L1D3PHI3Z2_L2D4PHI3Z1),
.stubpairout(TE_L1D3PHI3Z2_L2D4PHI3Z1_SP_L1D3PHI3Z2_L2D4PHI3Z1),
.valid_data(TE_L1D3PHI3Z2_L2D4PHI3Z1_SP_L1D3PHI3Z2_L2D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z2_L2D4PHI4Z1_phi.txt","TETable_TE_L1D3PHI3Z2_L2D4PHI4Z1_z.txt") TE_L1D3PHI3Z2_L2D4PHI4Z1(
.number_in1(VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1_number),
.read_add1(VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1_read_add),
.innervmstubin(VMS_L1D3PHI3Z2n4_TE_L1D3PHI3Z2_L2D4PHI4Z1),
.number_in2(VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1_number),
.read_add2(VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1_read_add),
.outervmstubin(VMS_L2D4PHI4Z1n2_TE_L1D3PHI3Z2_L2D4PHI4Z1),
.stubpairout(TE_L1D3PHI3Z2_L2D4PHI4Z1_SP_L1D3PHI3Z2_L2D4PHI4Z1),
.valid_data(TE_L1D3PHI3Z2_L2D4PHI4Z1_SP_L1D3PHI3Z2_L2D4PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z2_L2D4PHI1Z2_phi.txt","TETable_TE_L1D3PHI1Z2_L2D4PHI1Z2_z.txt") TE_L1D3PHI1Z2_L2D4PHI1Z2(
.number_in1(VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2_number),
.read_add1(VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2_read_add),
.innervmstubin(VMS_L1D3PHI1Z2n5_TE_L1D3PHI1Z2_L2D4PHI1Z2),
.number_in2(VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2_number),
.read_add2(VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2_read_add),
.outervmstubin(VMS_L2D4PHI1Z2n1_TE_L1D3PHI1Z2_L2D4PHI1Z2),
.stubpairout(TE_L1D3PHI1Z2_L2D4PHI1Z2_SP_L1D3PHI1Z2_L2D4PHI1Z2),
.valid_data(TE_L1D3PHI1Z2_L2D4PHI1Z2_SP_L1D3PHI1Z2_L2D4PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI1Z2_L2D4PHI2Z2_phi.txt","TETable_TE_L1D3PHI1Z2_L2D4PHI2Z2_z.txt") TE_L1D3PHI1Z2_L2D4PHI2Z2(
.number_in1(VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2_number),
.read_add1(VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2_read_add),
.innervmstubin(VMS_L1D3PHI1Z2n6_TE_L1D3PHI1Z2_L2D4PHI2Z2),
.number_in2(VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2_number),
.read_add2(VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2_read_add),
.outervmstubin(VMS_L2D4PHI2Z2n1_TE_L1D3PHI1Z2_L2D4PHI2Z2),
.stubpairout(TE_L1D3PHI1Z2_L2D4PHI2Z2_SP_L1D3PHI1Z2_L2D4PHI2Z2),
.valid_data(TE_L1D3PHI1Z2_L2D4PHI2Z2_SP_L1D3PHI1Z2_L2D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z2_L2D4PHI2Z2_phi.txt","TETable_TE_L1D3PHI2Z2_L2D4PHI2Z2_z.txt") TE_L1D3PHI2Z2_L2D4PHI2Z2(
.number_in1(VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2_number),
.read_add1(VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2_read_add),
.innervmstubin(VMS_L1D3PHI2Z2n5_TE_L1D3PHI2Z2_L2D4PHI2Z2),
.number_in2(VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2_number),
.read_add2(VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2_read_add),
.outervmstubin(VMS_L2D4PHI2Z2n2_TE_L1D3PHI2Z2_L2D4PHI2Z2),
.stubpairout(TE_L1D3PHI2Z2_L2D4PHI2Z2_SP_L1D3PHI2Z2_L2D4PHI2Z2),
.valid_data(TE_L1D3PHI2Z2_L2D4PHI2Z2_SP_L1D3PHI2Z2_L2D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI2Z2_L2D4PHI3Z2_phi.txt","TETable_TE_L1D3PHI2Z2_L2D4PHI3Z2_z.txt") TE_L1D3PHI2Z2_L2D4PHI3Z2(
.number_in1(VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2_number),
.read_add1(VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2_read_add),
.innervmstubin(VMS_L1D3PHI2Z2n6_TE_L1D3PHI2Z2_L2D4PHI3Z2),
.number_in2(VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2_number),
.read_add2(VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2_read_add),
.outervmstubin(VMS_L2D4PHI3Z2n1_TE_L1D3PHI2Z2_L2D4PHI3Z2),
.stubpairout(TE_L1D3PHI2Z2_L2D4PHI3Z2_SP_L1D3PHI2Z2_L2D4PHI3Z2),
.valid_data(TE_L1D3PHI2Z2_L2D4PHI3Z2_SP_L1D3PHI2Z2_L2D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z2_L2D4PHI3Z2_phi.txt","TETable_TE_L1D3PHI3Z2_L2D4PHI3Z2_z.txt") TE_L1D3PHI3Z2_L2D4PHI3Z2(
.number_in1(VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2_number),
.read_add1(VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2_read_add),
.innervmstubin(VMS_L1D3PHI3Z2n5_TE_L1D3PHI3Z2_L2D4PHI3Z2),
.number_in2(VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2_number),
.read_add2(VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2_read_add),
.outervmstubin(VMS_L2D4PHI3Z2n2_TE_L1D3PHI3Z2_L2D4PHI3Z2),
.stubpairout(TE_L1D3PHI3Z2_L2D4PHI3Z2_SP_L1D3PHI3Z2_L2D4PHI3Z2),
.valid_data(TE_L1D3PHI3Z2_L2D4PHI3Z2_SP_L1D3PHI3Z2_L2D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D3PHI3Z2_L2D4PHI4Z2_phi.txt","TETable_TE_L1D3PHI3Z2_L2D4PHI4Z2_z.txt") TE_L1D3PHI3Z2_L2D4PHI4Z2(
.number_in1(VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2_number),
.read_add1(VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2_read_add),
.innervmstubin(VMS_L1D3PHI3Z2n6_TE_L1D3PHI3Z2_L2D4PHI4Z2),
.number_in2(VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2_number),
.read_add2(VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2_read_add),
.outervmstubin(VMS_L2D4PHI4Z2n1_TE_L1D3PHI3Z2_L2D4PHI4Z2),
.stubpairout(TE_L1D3PHI3Z2_L2D4PHI4Z2_SP_L1D3PHI3Z2_L2D4PHI4Z2),
.valid_data(TE_L1D3PHI3Z2_L2D4PHI4Z2_SP_L1D3PHI3Z2_L2D4PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D4PHI1Z1_L2D4PHI1Z2_phi.txt","TETable_TE_L1D4PHI1Z1_L2D4PHI1Z2_z.txt") TE_L1D4PHI1Z1_L2D4PHI1Z2(
.number_in1(VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2_number),
.read_add1(VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2_read_add),
.outervmstubin(VMS_L2D4PHI1Z2n2_TE_L1D4PHI1Z1_L2D4PHI1Z2),
.number_in2(VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2_number),
.read_add2(VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2_read_add),
.innervmstubin(VMS_L1D4PHI1Z1n1_TE_L1D4PHI1Z1_L2D4PHI1Z2),
.stubpairout(TE_L1D4PHI1Z1_L2D4PHI1Z2_SP_L1D4PHI1Z1_L2D4PHI1Z2),
.valid_data(TE_L1D4PHI1Z1_L2D4PHI1Z2_SP_L1D4PHI1Z1_L2D4PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D4PHI1Z1_L2D4PHI2Z2_phi.txt","TETable_TE_L1D4PHI1Z1_L2D4PHI2Z2_z.txt") TE_L1D4PHI1Z1_L2D4PHI2Z2(
.number_in1(VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2_number),
.read_add1(VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2_read_add),
.outervmstubin(VMS_L2D4PHI2Z2n3_TE_L1D4PHI1Z1_L2D4PHI2Z2),
.number_in2(VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2_number),
.read_add2(VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2_read_add),
.innervmstubin(VMS_L1D4PHI1Z1n2_TE_L1D4PHI1Z1_L2D4PHI2Z2),
.stubpairout(TE_L1D4PHI1Z1_L2D4PHI2Z2_SP_L1D4PHI1Z1_L2D4PHI2Z2),
.valid_data(TE_L1D4PHI1Z1_L2D4PHI2Z2_SP_L1D4PHI1Z1_L2D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D4PHI2Z1_L2D4PHI2Z2_phi.txt","TETable_TE_L1D4PHI2Z1_L2D4PHI2Z2_z.txt") TE_L1D4PHI2Z1_L2D4PHI2Z2(
.number_in1(VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2_number),
.read_add1(VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2_read_add),
.outervmstubin(VMS_L2D4PHI2Z2n4_TE_L1D4PHI2Z1_L2D4PHI2Z2),
.number_in2(VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2_number),
.read_add2(VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2_read_add),
.innervmstubin(VMS_L1D4PHI2Z1n1_TE_L1D4PHI2Z1_L2D4PHI2Z2),
.stubpairout(TE_L1D4PHI2Z1_L2D4PHI2Z2_SP_L1D4PHI2Z1_L2D4PHI2Z2),
.valid_data(TE_L1D4PHI2Z1_L2D4PHI2Z2_SP_L1D4PHI2Z1_L2D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D4PHI2Z1_L2D4PHI3Z2_phi.txt","TETable_TE_L1D4PHI2Z1_L2D4PHI3Z2_z.txt") TE_L1D4PHI2Z1_L2D4PHI3Z2(
.number_in1(VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2_number),
.read_add1(VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2_read_add),
.outervmstubin(VMS_L2D4PHI3Z2n3_TE_L1D4PHI2Z1_L2D4PHI3Z2),
.number_in2(VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2_number),
.read_add2(VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2_read_add),
.innervmstubin(VMS_L1D4PHI2Z1n2_TE_L1D4PHI2Z1_L2D4PHI3Z2),
.stubpairout(TE_L1D4PHI2Z1_L2D4PHI3Z2_SP_L1D4PHI2Z1_L2D4PHI3Z2),
.valid_data(TE_L1D4PHI2Z1_L2D4PHI3Z2_SP_L1D4PHI2Z1_L2D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D4PHI3Z1_L2D4PHI3Z2_phi.txt","TETable_TE_L1D4PHI3Z1_L2D4PHI3Z2_z.txt") TE_L1D4PHI3Z1_L2D4PHI3Z2(
.number_in1(VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2_number),
.read_add1(VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2_read_add),
.outervmstubin(VMS_L2D4PHI3Z2n4_TE_L1D4PHI3Z1_L2D4PHI3Z2),
.number_in2(VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2_number),
.read_add2(VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2_read_add),
.innervmstubin(VMS_L1D4PHI3Z1n1_TE_L1D4PHI3Z1_L2D4PHI3Z2),
.stubpairout(TE_L1D4PHI3Z1_L2D4PHI3Z2_SP_L1D4PHI3Z1_L2D4PHI3Z2),
.valid_data(TE_L1D4PHI3Z1_L2D4PHI3Z2_SP_L1D4PHI3Z1_L2D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L1D4PHI3Z1_L2D4PHI4Z2_phi.txt","TETable_TE_L1D4PHI3Z1_L2D4PHI4Z2_z.txt") TE_L1D4PHI3Z1_L2D4PHI4Z2(
.number_in1(VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_number),
.read_add1(VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_read_add),
.outervmstubin(VMS_L2D4PHI4Z2n2_TE_L1D4PHI3Z1_L2D4PHI4Z2),
.number_in2(VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_number),
.read_add2(VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2_read_add),
.innervmstubin(VMS_L1D4PHI3Z1n2_TE_L1D4PHI3Z1_L2D4PHI4Z2),
.stubpairout(TE_L1D4PHI3Z1_L2D4PHI4Z2_SP_L1D4PHI3Z1_L2D4PHI4Z2),
.valid_data(TE_L1D4PHI3Z1_L2D4PHI4Z2_SP_L1D4PHI3Z1_L2D4PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI1Z1_L4D3PHI1Z1_phi.txt","TETable_TE_L3D3PHI1Z1_L4D3PHI1Z1_z.txt") TE_L3D3PHI1Z1_L4D3PHI1Z1(
.number_in1(VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_number),
.read_add1(VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_read_add),
.innervmstubin(VMS_L3D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1),
.number_in2(VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_number),
.read_add2(VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1_read_add),
.outervmstubin(VMS_L4D3PHI1Z1n1_TE_L3D3PHI1Z1_L4D3PHI1Z1),
.stubpairout(TE_L3D3PHI1Z1_L4D3PHI1Z1_SP_L3D3PHI1Z1_L4D3PHI1Z1),
.valid_data(TE_L3D3PHI1Z1_L4D3PHI1Z1_SP_L3D3PHI1Z1_L4D3PHI1Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI1Z1_L4D3PHI2Z1_phi.txt","TETable_TE_L3D3PHI1Z1_L4D3PHI2Z1_z.txt") TE_L3D3PHI1Z1_L4D3PHI2Z1(
.number_in1(VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1_number),
.read_add1(VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1_read_add),
.innervmstubin(VMS_L3D3PHI1Z1n2_TE_L3D3PHI1Z1_L4D3PHI2Z1),
.number_in2(VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1_number),
.read_add2(VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1_read_add),
.outervmstubin(VMS_L4D3PHI2Z1n1_TE_L3D3PHI1Z1_L4D3PHI2Z1),
.stubpairout(TE_L3D3PHI1Z1_L4D3PHI2Z1_SP_L3D3PHI1Z1_L4D3PHI2Z1),
.valid_data(TE_L3D3PHI1Z1_L4D3PHI2Z1_SP_L3D3PHI1Z1_L4D3PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI2Z1_L4D3PHI2Z1_phi.txt","TETable_TE_L3D3PHI2Z1_L4D3PHI2Z1_z.txt") TE_L3D3PHI2Z1_L4D3PHI2Z1(
.number_in1(VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1_number),
.read_add1(VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1_read_add),
.outervmstubin(VMS_L4D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI2Z1),
.number_in2(VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1_number),
.read_add2(VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1_read_add),
.innervmstubin(VMS_L3D3PHI2Z1n1_TE_L3D3PHI2Z1_L4D3PHI2Z1),
.stubpairout(TE_L3D3PHI2Z1_L4D3PHI2Z1_SP_L3D3PHI2Z1_L4D3PHI2Z1),
.valid_data(TE_L3D3PHI2Z1_L4D3PHI2Z1_SP_L3D3PHI2Z1_L4D3PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI2Z1_L4D3PHI3Z1_phi.txt","TETable_TE_L3D3PHI2Z1_L4D3PHI3Z1_z.txt") TE_L3D3PHI2Z1_L4D3PHI3Z1(
.number_in1(VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1_number),
.read_add1(VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1_read_add),
.innervmstubin(VMS_L3D3PHI2Z1n2_TE_L3D3PHI2Z1_L4D3PHI3Z1),
.number_in2(VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1_number),
.read_add2(VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1_read_add),
.outervmstubin(VMS_L4D3PHI3Z1n1_TE_L3D3PHI2Z1_L4D3PHI3Z1),
.stubpairout(TE_L3D3PHI2Z1_L4D3PHI3Z1_SP_L3D3PHI2Z1_L4D3PHI3Z1),
.valid_data(TE_L3D3PHI2Z1_L4D3PHI3Z1_SP_L3D3PHI2Z1_L4D3PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI3Z1_L4D3PHI3Z1_phi.txt","TETable_TE_L3D3PHI3Z1_L4D3PHI3Z1_z.txt") TE_L3D3PHI3Z1_L4D3PHI3Z1(
.number_in1(VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1_number),
.read_add1(VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1_read_add),
.outervmstubin(VMS_L4D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI3Z1),
.number_in2(VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1_number),
.read_add2(VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1_read_add),
.innervmstubin(VMS_L3D3PHI3Z1n1_TE_L3D3PHI3Z1_L4D3PHI3Z1),
.stubpairout(TE_L3D3PHI3Z1_L4D3PHI3Z1_SP_L3D3PHI3Z1_L4D3PHI3Z1),
.valid_data(TE_L3D3PHI3Z1_L4D3PHI3Z1_SP_L3D3PHI3Z1_L4D3PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI3Z1_L4D3PHI4Z1_phi.txt","TETable_TE_L3D3PHI3Z1_L4D3PHI4Z1_z.txt") TE_L3D3PHI3Z1_L4D3PHI4Z1(
.number_in1(VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1_number),
.read_add1(VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1_read_add),
.innervmstubin(VMS_L3D3PHI3Z1n2_TE_L3D3PHI3Z1_L4D3PHI4Z1),
.number_in2(VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1_number),
.read_add2(VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1_read_add),
.outervmstubin(VMS_L4D3PHI4Z1n1_TE_L3D3PHI3Z1_L4D3PHI4Z1),
.stubpairout(TE_L3D3PHI3Z1_L4D3PHI4Z1_SP_L3D3PHI3Z1_L4D3PHI4Z1),
.valid_data(TE_L3D3PHI3Z1_L4D3PHI4Z1_SP_L3D3PHI3Z1_L4D3PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI1Z2_L4D3PHI1Z2_phi.txt","TETable_TE_L3D3PHI1Z2_L4D3PHI1Z2_z.txt") TE_L3D3PHI1Z2_L4D3PHI1Z2(
.number_in1(VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_number),
.read_add1(VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_read_add),
.innervmstubin(VMS_L3D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2),
.number_in2(VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_number),
.read_add2(VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2_read_add),
.outervmstubin(VMS_L4D3PHI1Z2n1_TE_L3D3PHI1Z2_L4D3PHI1Z2),
.stubpairout(TE_L3D3PHI1Z2_L4D3PHI1Z2_SP_L3D3PHI1Z2_L4D3PHI1Z2),
.valid_data(TE_L3D3PHI1Z2_L4D3PHI1Z2_SP_L3D3PHI1Z2_L4D3PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI1Z2_L4D3PHI2Z2_phi.txt","TETable_TE_L3D3PHI1Z2_L4D3PHI2Z2_z.txt") TE_L3D3PHI1Z2_L4D3PHI2Z2(
.number_in1(VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2_number),
.read_add1(VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2_read_add),
.innervmstubin(VMS_L3D3PHI1Z2n2_TE_L3D3PHI1Z2_L4D3PHI2Z2),
.number_in2(VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2_number),
.read_add2(VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2_read_add),
.outervmstubin(VMS_L4D3PHI2Z2n1_TE_L3D3PHI1Z2_L4D3PHI2Z2),
.stubpairout(TE_L3D3PHI1Z2_L4D3PHI2Z2_SP_L3D3PHI1Z2_L4D3PHI2Z2),
.valid_data(TE_L3D3PHI1Z2_L4D3PHI2Z2_SP_L3D3PHI1Z2_L4D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI2Z2_L4D3PHI2Z2_phi.txt","TETable_TE_L3D3PHI2Z2_L4D3PHI2Z2_z.txt") TE_L3D3PHI2Z2_L4D3PHI2Z2(
.number_in1(VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2_number),
.read_add1(VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2_read_add),
.outervmstubin(VMS_L4D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI2Z2),
.number_in2(VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2_number),
.read_add2(VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2_read_add),
.innervmstubin(VMS_L3D3PHI2Z2n1_TE_L3D3PHI2Z2_L4D3PHI2Z2),
.stubpairout(TE_L3D3PHI2Z2_L4D3PHI2Z2_SP_L3D3PHI2Z2_L4D3PHI2Z2),
.valid_data(TE_L3D3PHI2Z2_L4D3PHI2Z2_SP_L3D3PHI2Z2_L4D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI2Z2_L4D3PHI3Z2_phi.txt","TETable_TE_L3D3PHI2Z2_L4D3PHI3Z2_z.txt") TE_L3D3PHI2Z2_L4D3PHI3Z2(
.number_in1(VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2_number),
.read_add1(VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2_read_add),
.innervmstubin(VMS_L3D3PHI2Z2n2_TE_L3D3PHI2Z2_L4D3PHI3Z2),
.number_in2(VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2_number),
.read_add2(VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2_read_add),
.outervmstubin(VMS_L4D3PHI3Z2n1_TE_L3D3PHI2Z2_L4D3PHI3Z2),
.stubpairout(TE_L3D3PHI2Z2_L4D3PHI3Z2_SP_L3D3PHI2Z2_L4D3PHI3Z2),
.valid_data(TE_L3D3PHI2Z2_L4D3PHI3Z2_SP_L3D3PHI2Z2_L4D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI3Z2_L4D3PHI3Z2_phi.txt","TETable_TE_L3D3PHI3Z2_L4D3PHI3Z2_z.txt") TE_L3D3PHI3Z2_L4D3PHI3Z2(
.number_in1(VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2_number),
.read_add1(VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2_read_add),
.outervmstubin(VMS_L4D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI3Z2),
.number_in2(VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2_number),
.read_add2(VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2_read_add),
.innervmstubin(VMS_L3D3PHI3Z2n1_TE_L3D3PHI3Z2_L4D3PHI3Z2),
.stubpairout(TE_L3D3PHI3Z2_L4D3PHI3Z2_SP_L3D3PHI3Z2_L4D3PHI3Z2),
.valid_data(TE_L3D3PHI3Z2_L4D3PHI3Z2_SP_L3D3PHI3Z2_L4D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI3Z2_L4D3PHI4Z2_phi.txt","TETable_TE_L3D3PHI3Z2_L4D3PHI4Z2_z.txt") TE_L3D3PHI3Z2_L4D3PHI4Z2(
.number_in1(VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2_number),
.read_add1(VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2_read_add),
.innervmstubin(VMS_L3D3PHI3Z2n2_TE_L3D3PHI3Z2_L4D3PHI4Z2),
.number_in2(VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2_number),
.read_add2(VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2_read_add),
.outervmstubin(VMS_L4D3PHI4Z2n1_TE_L3D3PHI3Z2_L4D3PHI4Z2),
.stubpairout(TE_L3D3PHI3Z2_L4D3PHI4Z2_SP_L3D3PHI3Z2_L4D3PHI4Z2),
.valid_data(TE_L3D3PHI3Z2_L4D3PHI4Z2_SP_L3D3PHI3Z2_L4D3PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI1Z1_L4D3PHI1Z2_phi.txt","TETable_TE_L3D3PHI1Z1_L4D3PHI1Z2_z.txt") TE_L3D3PHI1Z1_L4D3PHI1Z2(
.number_in1(VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2_number),
.read_add1(VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2_read_add),
.innervmstubin(VMS_L3D3PHI1Z1n3_TE_L3D3PHI1Z1_L4D3PHI1Z2),
.number_in2(VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2_number),
.read_add2(VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2_read_add),
.outervmstubin(VMS_L4D3PHI1Z2n2_TE_L3D3PHI1Z1_L4D3PHI1Z2),
.stubpairout(TE_L3D3PHI1Z1_L4D3PHI1Z2_SP_L3D3PHI1Z1_L4D3PHI1Z2),
.valid_data(TE_L3D3PHI1Z1_L4D3PHI1Z2_SP_L3D3PHI1Z1_L4D3PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI1Z1_L4D3PHI2Z2_phi.txt","TETable_TE_L3D3PHI1Z1_L4D3PHI2Z2_z.txt") TE_L3D3PHI1Z1_L4D3PHI2Z2(
.number_in1(VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2_number),
.read_add1(VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2_read_add),
.innervmstubin(VMS_L3D3PHI1Z1n4_TE_L3D3PHI1Z1_L4D3PHI2Z2),
.number_in2(VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2_number),
.read_add2(VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2_read_add),
.outervmstubin(VMS_L4D3PHI2Z2n3_TE_L3D3PHI1Z1_L4D3PHI2Z2),
.stubpairout(TE_L3D3PHI1Z1_L4D3PHI2Z2_SP_L3D3PHI1Z1_L4D3PHI2Z2),
.valid_data(TE_L3D3PHI1Z1_L4D3PHI2Z2_SP_L3D3PHI1Z1_L4D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI2Z1_L4D3PHI2Z2_phi.txt","TETable_TE_L3D3PHI2Z1_L4D3PHI2Z2_z.txt") TE_L3D3PHI2Z1_L4D3PHI2Z2(
.number_in1(VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2_number),
.read_add1(VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2_read_add),
.innervmstubin(VMS_L3D3PHI2Z1n3_TE_L3D3PHI2Z1_L4D3PHI2Z2),
.number_in2(VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2_number),
.read_add2(VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2_read_add),
.outervmstubin(VMS_L4D3PHI2Z2n4_TE_L3D3PHI2Z1_L4D3PHI2Z2),
.stubpairout(TE_L3D3PHI2Z1_L4D3PHI2Z2_SP_L3D3PHI2Z1_L4D3PHI2Z2),
.valid_data(TE_L3D3PHI2Z1_L4D3PHI2Z2_SP_L3D3PHI2Z1_L4D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI2Z1_L4D3PHI3Z2_phi.txt","TETable_TE_L3D3PHI2Z1_L4D3PHI3Z2_z.txt") TE_L3D3PHI2Z1_L4D3PHI3Z2(
.number_in1(VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2_number),
.read_add1(VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2_read_add),
.innervmstubin(VMS_L3D3PHI2Z1n4_TE_L3D3PHI2Z1_L4D3PHI3Z2),
.number_in2(VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2_number),
.read_add2(VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2_read_add),
.outervmstubin(VMS_L4D3PHI3Z2n3_TE_L3D3PHI2Z1_L4D3PHI3Z2),
.stubpairout(TE_L3D3PHI2Z1_L4D3PHI3Z2_SP_L3D3PHI2Z1_L4D3PHI3Z2),
.valid_data(TE_L3D3PHI2Z1_L4D3PHI3Z2_SP_L3D3PHI2Z1_L4D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI3Z1_L4D3PHI3Z2_phi.txt","TETable_TE_L3D3PHI3Z1_L4D3PHI3Z2_z.txt") TE_L3D3PHI3Z1_L4D3PHI3Z2(
.number_in1(VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2_number),
.read_add1(VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2_read_add),
.innervmstubin(VMS_L3D3PHI3Z1n3_TE_L3D3PHI3Z1_L4D3PHI3Z2),
.number_in2(VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2_number),
.read_add2(VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2_read_add),
.outervmstubin(VMS_L4D3PHI3Z2n4_TE_L3D3PHI3Z1_L4D3PHI3Z2),
.stubpairout(TE_L3D3PHI3Z1_L4D3PHI3Z2_SP_L3D3PHI3Z1_L4D3PHI3Z2),
.valid_data(TE_L3D3PHI3Z1_L4D3PHI3Z2_SP_L3D3PHI3Z1_L4D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI3Z1_L4D3PHI4Z2_phi.txt","TETable_TE_L3D3PHI3Z1_L4D3PHI4Z2_z.txt") TE_L3D3PHI3Z1_L4D3PHI4Z2(
.number_in1(VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2_number),
.read_add1(VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2_read_add),
.innervmstubin(VMS_L3D3PHI3Z1n4_TE_L3D3PHI3Z1_L4D3PHI4Z2),
.number_in2(VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2_number),
.read_add2(VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2_read_add),
.outervmstubin(VMS_L4D3PHI4Z2n2_TE_L3D3PHI3Z1_L4D3PHI4Z2),
.stubpairout(TE_L3D3PHI3Z1_L4D3PHI4Z2_SP_L3D3PHI3Z1_L4D3PHI4Z2),
.valid_data(TE_L3D3PHI3Z1_L4D3PHI4Z2_SP_L3D3PHI3Z1_L4D3PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI1Z2_L4D4PHI1Z1_phi.txt","TETable_TE_L3D3PHI1Z2_L4D4PHI1Z1_z.txt") TE_L3D3PHI1Z2_L4D4PHI1Z1(
.number_in1(VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1_number),
.read_add1(VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1_read_add),
.innervmstubin(VMS_L3D3PHI1Z2n3_TE_L3D3PHI1Z2_L4D4PHI1Z1),
.number_in2(VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1_number),
.read_add2(VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1_read_add),
.outervmstubin(VMS_L4D4PHI1Z1n1_TE_L3D3PHI1Z2_L4D4PHI1Z1),
.stubpairout(TE_L3D3PHI1Z2_L4D4PHI1Z1_SP_L3D3PHI1Z2_L4D4PHI1Z1),
.valid_data(TE_L3D3PHI1Z2_L4D4PHI1Z1_SP_L3D3PHI1Z2_L4D4PHI1Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI1Z2_L4D4PHI2Z1_phi.txt","TETable_TE_L3D3PHI1Z2_L4D4PHI2Z1_z.txt") TE_L3D3PHI1Z2_L4D4PHI2Z1(
.number_in1(VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1_number),
.read_add1(VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1_read_add),
.innervmstubin(VMS_L3D3PHI1Z2n4_TE_L3D3PHI1Z2_L4D4PHI2Z1),
.number_in2(VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1_number),
.read_add2(VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1_read_add),
.outervmstubin(VMS_L4D4PHI2Z1n1_TE_L3D3PHI1Z2_L4D4PHI2Z1),
.stubpairout(TE_L3D3PHI1Z2_L4D4PHI2Z1_SP_L3D3PHI1Z2_L4D4PHI2Z1),
.valid_data(TE_L3D3PHI1Z2_L4D4PHI2Z1_SP_L3D3PHI1Z2_L4D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI2Z2_L4D4PHI2Z1_phi.txt","TETable_TE_L3D3PHI2Z2_L4D4PHI2Z1_z.txt") TE_L3D3PHI2Z2_L4D4PHI2Z1(
.number_in1(VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1_number),
.read_add1(VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1_read_add),
.innervmstubin(VMS_L3D3PHI2Z2n3_TE_L3D3PHI2Z2_L4D4PHI2Z1),
.number_in2(VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1_number),
.read_add2(VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1_read_add),
.outervmstubin(VMS_L4D4PHI2Z1n2_TE_L3D3PHI2Z2_L4D4PHI2Z1),
.stubpairout(TE_L3D3PHI2Z2_L4D4PHI2Z1_SP_L3D3PHI2Z2_L4D4PHI2Z1),
.valid_data(TE_L3D3PHI2Z2_L4D4PHI2Z1_SP_L3D3PHI2Z2_L4D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI2Z2_L4D4PHI3Z1_phi.txt","TETable_TE_L3D3PHI2Z2_L4D4PHI3Z1_z.txt") TE_L3D3PHI2Z2_L4D4PHI3Z1(
.number_in1(VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1_number),
.read_add1(VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1_read_add),
.innervmstubin(VMS_L3D3PHI2Z2n4_TE_L3D3PHI2Z2_L4D4PHI3Z1),
.number_in2(VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1_number),
.read_add2(VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1_read_add),
.outervmstubin(VMS_L4D4PHI3Z1n1_TE_L3D3PHI2Z2_L4D4PHI3Z1),
.stubpairout(TE_L3D3PHI2Z2_L4D4PHI3Z1_SP_L3D3PHI2Z2_L4D4PHI3Z1),
.valid_data(TE_L3D3PHI2Z2_L4D4PHI3Z1_SP_L3D3PHI2Z2_L4D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI3Z2_L4D4PHI3Z1_phi.txt","TETable_TE_L3D3PHI3Z2_L4D4PHI3Z1_z.txt") TE_L3D3PHI3Z2_L4D4PHI3Z1(
.number_in1(VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1_number),
.read_add1(VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1_read_add),
.innervmstubin(VMS_L3D3PHI3Z2n3_TE_L3D3PHI3Z2_L4D4PHI3Z1),
.number_in2(VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1_number),
.read_add2(VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1_read_add),
.outervmstubin(VMS_L4D4PHI3Z1n2_TE_L3D3PHI3Z2_L4D4PHI3Z1),
.stubpairout(TE_L3D3PHI3Z2_L4D4PHI3Z1_SP_L3D3PHI3Z2_L4D4PHI3Z1),
.valid_data(TE_L3D3PHI3Z2_L4D4PHI3Z1_SP_L3D3PHI3Z2_L4D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D3PHI3Z2_L4D4PHI4Z1_phi.txt","TETable_TE_L3D3PHI3Z2_L4D4PHI4Z1_z.txt") TE_L3D3PHI3Z2_L4D4PHI4Z1(
.number_in1(VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1_number),
.read_add1(VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1_read_add),
.innervmstubin(VMS_L3D3PHI3Z2n4_TE_L3D3PHI3Z2_L4D4PHI4Z1),
.number_in2(VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1_number),
.read_add2(VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1_read_add),
.outervmstubin(VMS_L4D4PHI4Z1n1_TE_L3D3PHI3Z2_L4D4PHI4Z1),
.stubpairout(TE_L3D3PHI3Z2_L4D4PHI4Z1_SP_L3D3PHI3Z2_L4D4PHI4Z1),
.valid_data(TE_L3D3PHI3Z2_L4D4PHI4Z1_SP_L3D3PHI3Z2_L4D4PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI1Z1_L4D4PHI1Z1_phi.txt","TETable_TE_L3D4PHI1Z1_L4D4PHI1Z1_z.txt") TE_L3D4PHI1Z1_L4D4PHI1Z1(
.number_in1(VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1_number),
.read_add1(VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1_read_add),
.outervmstubin(VMS_L4D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI1Z1),
.number_in2(VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1_number),
.read_add2(VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1_read_add),
.innervmstubin(VMS_L3D4PHI1Z1n1_TE_L3D4PHI1Z1_L4D4PHI1Z1),
.stubpairout(TE_L3D4PHI1Z1_L4D4PHI1Z1_SP_L3D4PHI1Z1_L4D4PHI1Z1),
.valid_data(TE_L3D4PHI1Z1_L4D4PHI1Z1_SP_L3D4PHI1Z1_L4D4PHI1Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI1Z1_L4D4PHI2Z1_phi.txt","TETable_TE_L3D4PHI1Z1_L4D4PHI2Z1_z.txt") TE_L3D4PHI1Z1_L4D4PHI2Z1(
.number_in1(VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1_number),
.read_add1(VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1_read_add),
.outervmstubin(VMS_L4D4PHI2Z1n3_TE_L3D4PHI1Z1_L4D4PHI2Z1),
.number_in2(VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1_number),
.read_add2(VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1_read_add),
.innervmstubin(VMS_L3D4PHI1Z1n2_TE_L3D4PHI1Z1_L4D4PHI2Z1),
.stubpairout(TE_L3D4PHI1Z1_L4D4PHI2Z1_SP_L3D4PHI1Z1_L4D4PHI2Z1),
.valid_data(TE_L3D4PHI1Z1_L4D4PHI2Z1_SP_L3D4PHI1Z1_L4D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI2Z1_L4D4PHI2Z1_phi.txt","TETable_TE_L3D4PHI2Z1_L4D4PHI2Z1_z.txt") TE_L3D4PHI2Z1_L4D4PHI2Z1(
.number_in1(VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1_number),
.read_add1(VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1_read_add),
.outervmstubin(VMS_L4D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI2Z1),
.number_in2(VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1_number),
.read_add2(VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1_read_add),
.innervmstubin(VMS_L3D4PHI2Z1n1_TE_L3D4PHI2Z1_L4D4PHI2Z1),
.stubpairout(TE_L3D4PHI2Z1_L4D4PHI2Z1_SP_L3D4PHI2Z1_L4D4PHI2Z1),
.valid_data(TE_L3D4PHI2Z1_L4D4PHI2Z1_SP_L3D4PHI2Z1_L4D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI2Z1_L4D4PHI3Z1_phi.txt","TETable_TE_L3D4PHI2Z1_L4D4PHI3Z1_z.txt") TE_L3D4PHI2Z1_L4D4PHI3Z1(
.number_in1(VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1_number),
.read_add1(VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1_read_add),
.outervmstubin(VMS_L4D4PHI3Z1n3_TE_L3D4PHI2Z1_L4D4PHI3Z1),
.number_in2(VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1_number),
.read_add2(VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1_read_add),
.innervmstubin(VMS_L3D4PHI2Z1n2_TE_L3D4PHI2Z1_L4D4PHI3Z1),
.stubpairout(TE_L3D4PHI2Z1_L4D4PHI3Z1_SP_L3D4PHI2Z1_L4D4PHI3Z1),
.valid_data(TE_L3D4PHI2Z1_L4D4PHI3Z1_SP_L3D4PHI2Z1_L4D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI3Z1_L4D4PHI3Z1_phi.txt","TETable_TE_L3D4PHI3Z1_L4D4PHI3Z1_z.txt") TE_L3D4PHI3Z1_L4D4PHI3Z1(
.number_in1(VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1_number),
.read_add1(VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1_read_add),
.outervmstubin(VMS_L4D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI3Z1),
.number_in2(VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1_number),
.read_add2(VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1_read_add),
.innervmstubin(VMS_L3D4PHI3Z1n1_TE_L3D4PHI3Z1_L4D4PHI3Z1),
.stubpairout(TE_L3D4PHI3Z1_L4D4PHI3Z1_SP_L3D4PHI3Z1_L4D4PHI3Z1),
.valid_data(TE_L3D4PHI3Z1_L4D4PHI3Z1_SP_L3D4PHI3Z1_L4D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI3Z1_L4D4PHI4Z1_phi.txt","TETable_TE_L3D4PHI3Z1_L4D4PHI4Z1_z.txt") TE_L3D4PHI3Z1_L4D4PHI4Z1(
.number_in1(VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_number),
.read_add1(VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_read_add),
.outervmstubin(VMS_L4D4PHI4Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1),
.number_in2(VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_number),
.read_add2(VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1_read_add),
.innervmstubin(VMS_L3D4PHI3Z1n2_TE_L3D4PHI3Z1_L4D4PHI4Z1),
.stubpairout(TE_L3D4PHI3Z1_L4D4PHI4Z1_SP_L3D4PHI3Z1_L4D4PHI4Z1),
.valid_data(TE_L3D4PHI3Z1_L4D4PHI4Z1_SP_L3D4PHI3Z1_L4D4PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI1Z1_L4D4PHI1Z2_phi.txt","TETable_TE_L3D4PHI1Z1_L4D4PHI1Z2_z.txt") TE_L3D4PHI1Z1_L4D4PHI1Z2(
.number_in1(VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2_number),
.read_add1(VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2_read_add),
.innervmstubin(VMS_L3D4PHI1Z1n3_TE_L3D4PHI1Z1_L4D4PHI1Z2),
.number_in2(VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2_number),
.read_add2(VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2_read_add),
.outervmstubin(VMS_L4D4PHI1Z2n1_TE_L3D4PHI1Z1_L4D4PHI1Z2),
.stubpairout(TE_L3D4PHI1Z1_L4D4PHI1Z2_SP_L3D4PHI1Z1_L4D4PHI1Z2),
.valid_data(TE_L3D4PHI1Z1_L4D4PHI1Z2_SP_L3D4PHI1Z1_L4D4PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI1Z1_L4D4PHI2Z2_phi.txt","TETable_TE_L3D4PHI1Z1_L4D4PHI2Z2_z.txt") TE_L3D4PHI1Z1_L4D4PHI2Z2(
.number_in1(VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2_number),
.read_add1(VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2_read_add),
.innervmstubin(VMS_L3D4PHI1Z1n4_TE_L3D4PHI1Z1_L4D4PHI2Z2),
.number_in2(VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2_number),
.read_add2(VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2_read_add),
.outervmstubin(VMS_L4D4PHI2Z2n1_TE_L3D4PHI1Z1_L4D4PHI2Z2),
.stubpairout(TE_L3D4PHI1Z1_L4D4PHI2Z2_SP_L3D4PHI1Z1_L4D4PHI2Z2),
.valid_data(TE_L3D4PHI1Z1_L4D4PHI2Z2_SP_L3D4PHI1Z1_L4D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI2Z1_L4D4PHI2Z2_phi.txt","TETable_TE_L3D4PHI2Z1_L4D4PHI2Z2_z.txt") TE_L3D4PHI2Z1_L4D4PHI2Z2(
.number_in1(VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2_number),
.read_add1(VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2_read_add),
.innervmstubin(VMS_L3D4PHI2Z1n3_TE_L3D4PHI2Z1_L4D4PHI2Z2),
.number_in2(VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2_number),
.read_add2(VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2_read_add),
.outervmstubin(VMS_L4D4PHI2Z2n2_TE_L3D4PHI2Z1_L4D4PHI2Z2),
.stubpairout(TE_L3D4PHI2Z1_L4D4PHI2Z2_SP_L3D4PHI2Z1_L4D4PHI2Z2),
.valid_data(TE_L3D4PHI2Z1_L4D4PHI2Z2_SP_L3D4PHI2Z1_L4D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI2Z1_L4D4PHI3Z2_phi.txt","TETable_TE_L3D4PHI2Z1_L4D4PHI3Z2_z.txt") TE_L3D4PHI2Z1_L4D4PHI3Z2(
.number_in1(VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2_number),
.read_add1(VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2_read_add),
.innervmstubin(VMS_L3D4PHI2Z1n4_TE_L3D4PHI2Z1_L4D4PHI3Z2),
.number_in2(VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2_number),
.read_add2(VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2_read_add),
.outervmstubin(VMS_L4D4PHI3Z2n1_TE_L3D4PHI2Z1_L4D4PHI3Z2),
.stubpairout(TE_L3D4PHI2Z1_L4D4PHI3Z2_SP_L3D4PHI2Z1_L4D4PHI3Z2),
.valid_data(TE_L3D4PHI2Z1_L4D4PHI3Z2_SP_L3D4PHI2Z1_L4D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI3Z1_L4D4PHI3Z2_phi.txt","TETable_TE_L3D4PHI3Z1_L4D4PHI3Z2_z.txt") TE_L3D4PHI3Z1_L4D4PHI3Z2(
.number_in1(VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2_number),
.read_add1(VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2_read_add),
.innervmstubin(VMS_L3D4PHI3Z1n3_TE_L3D4PHI3Z1_L4D4PHI3Z2),
.number_in2(VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2_number),
.read_add2(VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2_read_add),
.outervmstubin(VMS_L4D4PHI3Z2n2_TE_L3D4PHI3Z1_L4D4PHI3Z2),
.stubpairout(TE_L3D4PHI3Z1_L4D4PHI3Z2_SP_L3D4PHI3Z1_L4D4PHI3Z2),
.valid_data(TE_L3D4PHI3Z1_L4D4PHI3Z2_SP_L3D4PHI3Z1_L4D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI3Z1_L4D4PHI4Z2_phi.txt","TETable_TE_L3D4PHI3Z1_L4D4PHI4Z2_z.txt") TE_L3D4PHI3Z1_L4D4PHI4Z2(
.number_in1(VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2_number),
.read_add1(VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2_read_add),
.innervmstubin(VMS_L3D4PHI3Z1n4_TE_L3D4PHI3Z1_L4D4PHI4Z2),
.number_in2(VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2_number),
.read_add2(VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2_read_add),
.outervmstubin(VMS_L4D4PHI4Z2n1_TE_L3D4PHI3Z1_L4D4PHI4Z2),
.stubpairout(TE_L3D4PHI3Z1_L4D4PHI4Z2_SP_L3D4PHI3Z1_L4D4PHI4Z2),
.valid_data(TE_L3D4PHI3Z1_L4D4PHI4Z2_SP_L3D4PHI3Z1_L4D4PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI1Z2_L4D4PHI1Z2_phi.txt","TETable_TE_L3D4PHI1Z2_L4D4PHI1Z2_z.txt") TE_L3D4PHI1Z2_L4D4PHI1Z2(
.number_in1(VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2_number),
.read_add1(VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2_read_add),
.outervmstubin(VMS_L4D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI1Z2),
.number_in2(VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2_number),
.read_add2(VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2_read_add),
.innervmstubin(VMS_L3D4PHI1Z2n1_TE_L3D4PHI1Z2_L4D4PHI1Z2),
.stubpairout(TE_L3D4PHI1Z2_L4D4PHI1Z2_SP_L3D4PHI1Z2_L4D4PHI1Z2),
.valid_data(TE_L3D4PHI1Z2_L4D4PHI1Z2_SP_L3D4PHI1Z2_L4D4PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI1Z2_L4D4PHI2Z2_phi.txt","TETable_TE_L3D4PHI1Z2_L4D4PHI2Z2_z.txt") TE_L3D4PHI1Z2_L4D4PHI2Z2(
.number_in1(VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2_number),
.read_add1(VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2_read_add),
.outervmstubin(VMS_L4D4PHI2Z2n3_TE_L3D4PHI1Z2_L4D4PHI2Z2),
.number_in2(VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2_number),
.read_add2(VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2_read_add),
.innervmstubin(VMS_L3D4PHI1Z2n2_TE_L3D4PHI1Z2_L4D4PHI2Z2),
.stubpairout(TE_L3D4PHI1Z2_L4D4PHI2Z2_SP_L3D4PHI1Z2_L4D4PHI2Z2),
.valid_data(TE_L3D4PHI1Z2_L4D4PHI2Z2_SP_L3D4PHI1Z2_L4D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI2Z2_L4D4PHI2Z2_phi.txt","TETable_TE_L3D4PHI2Z2_L4D4PHI2Z2_z.txt") TE_L3D4PHI2Z2_L4D4PHI2Z2(
.number_in1(VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2_number),
.read_add1(VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2_read_add),
.outervmstubin(VMS_L4D4PHI2Z2n4_TE_L3D4PHI2Z2_L4D4PHI2Z2),
.number_in2(VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2_number),
.read_add2(VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2_read_add),
.innervmstubin(VMS_L3D4PHI2Z2n1_TE_L3D4PHI2Z2_L4D4PHI2Z2),
.stubpairout(TE_L3D4PHI2Z2_L4D4PHI2Z2_SP_L3D4PHI2Z2_L4D4PHI2Z2),
.valid_data(TE_L3D4PHI2Z2_L4D4PHI2Z2_SP_L3D4PHI2Z2_L4D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI2Z2_L4D4PHI3Z2_phi.txt","TETable_TE_L3D4PHI2Z2_L4D4PHI3Z2_z.txt") TE_L3D4PHI2Z2_L4D4PHI3Z2(
.number_in1(VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2_number),
.read_add1(VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2_read_add),
.outervmstubin(VMS_L4D4PHI3Z2n3_TE_L3D4PHI2Z2_L4D4PHI3Z2),
.number_in2(VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2_number),
.read_add2(VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2_read_add),
.innervmstubin(VMS_L3D4PHI2Z2n2_TE_L3D4PHI2Z2_L4D4PHI3Z2),
.stubpairout(TE_L3D4PHI2Z2_L4D4PHI3Z2_SP_L3D4PHI2Z2_L4D4PHI3Z2),
.valid_data(TE_L3D4PHI2Z2_L4D4PHI3Z2_SP_L3D4PHI2Z2_L4D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI3Z2_L4D4PHI3Z2_phi.txt","TETable_TE_L3D4PHI3Z2_L4D4PHI3Z2_z.txt") TE_L3D4PHI3Z2_L4D4PHI3Z2(
.number_in1(VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2_number),
.read_add1(VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2_read_add),
.outervmstubin(VMS_L4D4PHI3Z2n4_TE_L3D4PHI3Z2_L4D4PHI3Z2),
.number_in2(VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2_number),
.read_add2(VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2_read_add),
.innervmstubin(VMS_L3D4PHI3Z2n1_TE_L3D4PHI3Z2_L4D4PHI3Z2),
.stubpairout(TE_L3D4PHI3Z2_L4D4PHI3Z2_SP_L3D4PHI3Z2_L4D4PHI3Z2),
.valid_data(TE_L3D4PHI3Z2_L4D4PHI3Z2_SP_L3D4PHI3Z2_L4D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L3D4PHI3Z2_L4D4PHI4Z2_phi.txt","TETable_TE_L3D4PHI3Z2_L4D4PHI4Z2_z.txt") TE_L3D4PHI3Z2_L4D4PHI4Z2(
.number_in1(VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_number),
.read_add1(VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_read_add),
.outervmstubin(VMS_L4D4PHI4Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2),
.number_in2(VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_number),
.read_add2(VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2_read_add),
.innervmstubin(VMS_L3D4PHI3Z2n2_TE_L3D4PHI3Z2_L4D4PHI4Z2),
.stubpairout(TE_L3D4PHI3Z2_L4D4PHI4Z2_SP_L3D4PHI3Z2_L4D4PHI4Z2),
.valid_data(TE_L3D4PHI3Z2_L4D4PHI4Z2_SP_L3D4PHI3Z2_L4D4PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI1Z1_L6D3PHI1Z1_phi.txt","TETable_TE_L5D3PHI1Z1_L6D3PHI1Z1_z.txt") TE_L5D3PHI1Z1_L6D3PHI1Z1(
.number_in1(VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_number),
.read_add1(VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_read_add),
.innervmstubin(VMS_L5D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1),
.number_in2(VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_number),
.read_add2(VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1_read_add),
.outervmstubin(VMS_L6D3PHI1Z1n1_TE_L5D3PHI1Z1_L6D3PHI1Z1),
.stubpairout(TE_L5D3PHI1Z1_L6D3PHI1Z1_SP_L5D3PHI1Z1_L6D3PHI1Z1),
.valid_data(TE_L5D3PHI1Z1_L6D3PHI1Z1_SP_L5D3PHI1Z1_L6D3PHI1Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI1Z1_L6D3PHI2Z1_phi.txt","TETable_TE_L5D3PHI1Z1_L6D3PHI2Z1_z.txt") TE_L5D3PHI1Z1_L6D3PHI2Z1(
.number_in1(VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1_number),
.read_add1(VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1_read_add),
.innervmstubin(VMS_L5D3PHI1Z1n2_TE_L5D3PHI1Z1_L6D3PHI2Z1),
.number_in2(VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1_number),
.read_add2(VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1_read_add),
.outervmstubin(VMS_L6D3PHI2Z1n1_TE_L5D3PHI1Z1_L6D3PHI2Z1),
.stubpairout(TE_L5D3PHI1Z1_L6D3PHI2Z1_SP_L5D3PHI1Z1_L6D3PHI2Z1),
.valid_data(TE_L5D3PHI1Z1_L6D3PHI2Z1_SP_L5D3PHI1Z1_L6D3PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI2Z1_L6D3PHI2Z1_phi.txt","TETable_TE_L5D3PHI2Z1_L6D3PHI2Z1_z.txt") TE_L5D3PHI2Z1_L6D3PHI2Z1(
.number_in1(VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1_number),
.read_add1(VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1_read_add),
.outervmstubin(VMS_L6D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI2Z1),
.number_in2(VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1_number),
.read_add2(VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1_read_add),
.innervmstubin(VMS_L5D3PHI2Z1n1_TE_L5D3PHI2Z1_L6D3PHI2Z1),
.stubpairout(TE_L5D3PHI2Z1_L6D3PHI2Z1_SP_L5D3PHI2Z1_L6D3PHI2Z1),
.valid_data(TE_L5D3PHI2Z1_L6D3PHI2Z1_SP_L5D3PHI2Z1_L6D3PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI2Z1_L6D3PHI3Z1_phi.txt","TETable_TE_L5D3PHI2Z1_L6D3PHI3Z1_z.txt") TE_L5D3PHI2Z1_L6D3PHI3Z1(
.number_in1(VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1_number),
.read_add1(VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1_read_add),
.innervmstubin(VMS_L5D3PHI2Z1n2_TE_L5D3PHI2Z1_L6D3PHI3Z1),
.number_in2(VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1_number),
.read_add2(VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1_read_add),
.outervmstubin(VMS_L6D3PHI3Z1n1_TE_L5D3PHI2Z1_L6D3PHI3Z1),
.stubpairout(TE_L5D3PHI2Z1_L6D3PHI3Z1_SP_L5D3PHI2Z1_L6D3PHI3Z1),
.valid_data(TE_L5D3PHI2Z1_L6D3PHI3Z1_SP_L5D3PHI2Z1_L6D3PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI3Z1_L6D3PHI3Z1_phi.txt","TETable_TE_L5D3PHI3Z1_L6D3PHI3Z1_z.txt") TE_L5D3PHI3Z1_L6D3PHI3Z1(
.number_in1(VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1_number),
.read_add1(VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1_read_add),
.outervmstubin(VMS_L6D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI3Z1),
.number_in2(VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1_number),
.read_add2(VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1_read_add),
.innervmstubin(VMS_L5D3PHI3Z1n1_TE_L5D3PHI3Z1_L6D3PHI3Z1),
.stubpairout(TE_L5D3PHI3Z1_L6D3PHI3Z1_SP_L5D3PHI3Z1_L6D3PHI3Z1),
.valid_data(TE_L5D3PHI3Z1_L6D3PHI3Z1_SP_L5D3PHI3Z1_L6D3PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI3Z1_L6D3PHI4Z1_phi.txt","TETable_TE_L5D3PHI3Z1_L6D3PHI4Z1_z.txt") TE_L5D3PHI3Z1_L6D3PHI4Z1(
.number_in1(VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1_number),
.read_add1(VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1_read_add),
.innervmstubin(VMS_L5D3PHI3Z1n2_TE_L5D3PHI3Z1_L6D3PHI4Z1),
.number_in2(VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1_number),
.read_add2(VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1_read_add),
.outervmstubin(VMS_L6D3PHI4Z1n1_TE_L5D3PHI3Z1_L6D3PHI4Z1),
.stubpairout(TE_L5D3PHI3Z1_L6D3PHI4Z1_SP_L5D3PHI3Z1_L6D3PHI4Z1),
.valid_data(TE_L5D3PHI3Z1_L6D3PHI4Z1_SP_L5D3PHI3Z1_L6D3PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI1Z1_L6D3PHI1Z2_phi.txt","TETable_TE_L5D3PHI1Z1_L6D3PHI1Z2_z.txt") TE_L5D3PHI1Z1_L6D3PHI1Z2(
.number_in1(VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2_number),
.read_add1(VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2_read_add),
.innervmstubin(VMS_L5D3PHI1Z1n3_TE_L5D3PHI1Z1_L6D3PHI1Z2),
.number_in2(VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2_number),
.read_add2(VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2_read_add),
.outervmstubin(VMS_L6D3PHI1Z2n1_TE_L5D3PHI1Z1_L6D3PHI1Z2),
.stubpairout(TE_L5D3PHI1Z1_L6D3PHI1Z2_SP_L5D3PHI1Z1_L6D3PHI1Z2),
.valid_data(TE_L5D3PHI1Z1_L6D3PHI1Z2_SP_L5D3PHI1Z1_L6D3PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI1Z1_L6D3PHI2Z2_phi.txt","TETable_TE_L5D3PHI1Z1_L6D3PHI2Z2_z.txt") TE_L5D3PHI1Z1_L6D3PHI2Z2(
.number_in1(VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2_number),
.read_add1(VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2_read_add),
.innervmstubin(VMS_L5D3PHI1Z1n4_TE_L5D3PHI1Z1_L6D3PHI2Z2),
.number_in2(VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2_number),
.read_add2(VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2_read_add),
.outervmstubin(VMS_L6D3PHI2Z2n1_TE_L5D3PHI1Z1_L6D3PHI2Z2),
.stubpairout(TE_L5D3PHI1Z1_L6D3PHI2Z2_SP_L5D3PHI1Z1_L6D3PHI2Z2),
.valid_data(TE_L5D3PHI1Z1_L6D3PHI2Z2_SP_L5D3PHI1Z1_L6D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI2Z1_L6D3PHI2Z2_phi.txt","TETable_TE_L5D3PHI2Z1_L6D3PHI2Z2_z.txt") TE_L5D3PHI2Z1_L6D3PHI2Z2(
.number_in1(VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2_number),
.read_add1(VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2_read_add),
.innervmstubin(VMS_L5D3PHI2Z1n3_TE_L5D3PHI2Z1_L6D3PHI2Z2),
.number_in2(VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2_number),
.read_add2(VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2_read_add),
.outervmstubin(VMS_L6D3PHI2Z2n2_TE_L5D3PHI2Z1_L6D3PHI2Z2),
.stubpairout(TE_L5D3PHI2Z1_L6D3PHI2Z2_SP_L5D3PHI2Z1_L6D3PHI2Z2),
.valid_data(TE_L5D3PHI2Z1_L6D3PHI2Z2_SP_L5D3PHI2Z1_L6D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI2Z1_L6D3PHI3Z2_phi.txt","TETable_TE_L5D3PHI2Z1_L6D3PHI3Z2_z.txt") TE_L5D3PHI2Z1_L6D3PHI3Z2(
.number_in1(VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2_number),
.read_add1(VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2_read_add),
.innervmstubin(VMS_L5D3PHI2Z1n4_TE_L5D3PHI2Z1_L6D3PHI3Z2),
.number_in2(VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2_number),
.read_add2(VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2_read_add),
.outervmstubin(VMS_L6D3PHI3Z2n1_TE_L5D3PHI2Z1_L6D3PHI3Z2),
.stubpairout(TE_L5D3PHI2Z1_L6D3PHI3Z2_SP_L5D3PHI2Z1_L6D3PHI3Z2),
.valid_data(TE_L5D3PHI2Z1_L6D3PHI3Z2_SP_L5D3PHI2Z1_L6D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI3Z1_L6D3PHI3Z2_phi.txt","TETable_TE_L5D3PHI3Z1_L6D3PHI3Z2_z.txt") TE_L5D3PHI3Z1_L6D3PHI3Z2(
.number_in1(VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2_number),
.read_add1(VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2_read_add),
.innervmstubin(VMS_L5D3PHI3Z1n3_TE_L5D3PHI3Z1_L6D3PHI3Z2),
.number_in2(VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2_number),
.read_add2(VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2_read_add),
.outervmstubin(VMS_L6D3PHI3Z2n2_TE_L5D3PHI3Z1_L6D3PHI3Z2),
.stubpairout(TE_L5D3PHI3Z1_L6D3PHI3Z2_SP_L5D3PHI3Z1_L6D3PHI3Z2),
.valid_data(TE_L5D3PHI3Z1_L6D3PHI3Z2_SP_L5D3PHI3Z1_L6D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI3Z1_L6D3PHI4Z2_phi.txt","TETable_TE_L5D3PHI3Z1_L6D3PHI4Z2_z.txt") TE_L5D3PHI3Z1_L6D3PHI4Z2(
.number_in1(VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2_number),
.read_add1(VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2_read_add),
.innervmstubin(VMS_L5D3PHI3Z1n4_TE_L5D3PHI3Z1_L6D3PHI4Z2),
.number_in2(VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2_number),
.read_add2(VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2_read_add),
.outervmstubin(VMS_L6D3PHI4Z2n1_TE_L5D3PHI3Z1_L6D3PHI4Z2),
.stubpairout(TE_L5D3PHI3Z1_L6D3PHI4Z2_SP_L5D3PHI3Z1_L6D3PHI4Z2),
.valid_data(TE_L5D3PHI3Z1_L6D3PHI4Z2_SP_L5D3PHI3Z1_L6D3PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI1Z2_L6D3PHI1Z2_phi.txt","TETable_TE_L5D3PHI1Z2_L6D3PHI1Z2_z.txt") TE_L5D3PHI1Z2_L6D3PHI1Z2(
.number_in1(VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2_number),
.read_add1(VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2_read_add),
.outervmstubin(VMS_L6D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI1Z2),
.number_in2(VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2_number),
.read_add2(VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2_read_add),
.innervmstubin(VMS_L5D3PHI1Z2n1_TE_L5D3PHI1Z2_L6D3PHI1Z2),
.stubpairout(TE_L5D3PHI1Z2_L6D3PHI1Z2_SP_L5D3PHI1Z2_L6D3PHI1Z2),
.valid_data(TE_L5D3PHI1Z2_L6D3PHI1Z2_SP_L5D3PHI1Z2_L6D3PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI1Z2_L6D3PHI2Z2_phi.txt","TETable_TE_L5D3PHI1Z2_L6D3PHI2Z2_z.txt") TE_L5D3PHI1Z2_L6D3PHI2Z2(
.number_in1(VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2_number),
.read_add1(VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2_read_add),
.outervmstubin(VMS_L6D3PHI2Z2n3_TE_L5D3PHI1Z2_L6D3PHI2Z2),
.number_in2(VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2_number),
.read_add2(VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2_read_add),
.innervmstubin(VMS_L5D3PHI1Z2n2_TE_L5D3PHI1Z2_L6D3PHI2Z2),
.stubpairout(TE_L5D3PHI1Z2_L6D3PHI2Z2_SP_L5D3PHI1Z2_L6D3PHI2Z2),
.valid_data(TE_L5D3PHI1Z2_L6D3PHI2Z2_SP_L5D3PHI1Z2_L6D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI2Z2_L6D3PHI2Z2_phi.txt","TETable_TE_L5D3PHI2Z2_L6D3PHI2Z2_z.txt") TE_L5D3PHI2Z2_L6D3PHI2Z2(
.number_in1(VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2_number),
.read_add1(VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2_read_add),
.outervmstubin(VMS_L6D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D3PHI2Z2),
.number_in2(VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2_number),
.read_add2(VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2_read_add),
.innervmstubin(VMS_L5D3PHI2Z2n1_TE_L5D3PHI2Z2_L6D3PHI2Z2),
.stubpairout(TE_L5D3PHI2Z2_L6D3PHI2Z2_SP_L5D3PHI2Z2_L6D3PHI2Z2),
.valid_data(TE_L5D3PHI2Z2_L6D3PHI2Z2_SP_L5D3PHI2Z2_L6D3PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI2Z2_L6D3PHI3Z2_phi.txt","TETable_TE_L5D3PHI2Z2_L6D3PHI3Z2_z.txt") TE_L5D3PHI2Z2_L6D3PHI3Z2(
.number_in1(VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2_number),
.read_add1(VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2_read_add),
.outervmstubin(VMS_L6D3PHI3Z2n3_TE_L5D3PHI2Z2_L6D3PHI3Z2),
.number_in2(VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2_number),
.read_add2(VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2_read_add),
.innervmstubin(VMS_L5D3PHI2Z2n2_TE_L5D3PHI2Z2_L6D3PHI3Z2),
.stubpairout(TE_L5D3PHI2Z2_L6D3PHI3Z2_SP_L5D3PHI2Z2_L6D3PHI3Z2),
.valid_data(TE_L5D3PHI2Z2_L6D3PHI3Z2_SP_L5D3PHI2Z2_L6D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI3Z2_L6D3PHI3Z2_phi.txt","TETable_TE_L5D3PHI3Z2_L6D3PHI3Z2_z.txt") TE_L5D3PHI3Z2_L6D3PHI3Z2(
.number_in1(VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2_number),
.read_add1(VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2_read_add),
.outervmstubin(VMS_L6D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D3PHI3Z2),
.number_in2(VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2_number),
.read_add2(VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2_read_add),
.innervmstubin(VMS_L5D3PHI3Z2n1_TE_L5D3PHI3Z2_L6D3PHI3Z2),
.stubpairout(TE_L5D3PHI3Z2_L6D3PHI3Z2_SP_L5D3PHI3Z2_L6D3PHI3Z2),
.valid_data(TE_L5D3PHI3Z2_L6D3PHI3Z2_SP_L5D3PHI3Z2_L6D3PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI3Z2_L6D3PHI4Z2_phi.txt","TETable_TE_L5D3PHI3Z2_L6D3PHI4Z2_z.txt") TE_L5D3PHI3Z2_L6D3PHI4Z2(
.number_in1(VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_number),
.read_add1(VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_read_add),
.outervmstubin(VMS_L6D3PHI4Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2),
.number_in2(VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_number),
.read_add2(VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2_read_add),
.innervmstubin(VMS_L5D3PHI3Z2n2_TE_L5D3PHI3Z2_L6D3PHI4Z2),
.stubpairout(TE_L5D3PHI3Z2_L6D3PHI4Z2_SP_L5D3PHI3Z2_L6D3PHI4Z2),
.valid_data(TE_L5D3PHI3Z2_L6D3PHI4Z2_SP_L5D3PHI3Z2_L6D3PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI1Z2_L6D4PHI1Z1_phi.txt","TETable_TE_L5D3PHI1Z2_L6D4PHI1Z1_z.txt") TE_L5D3PHI1Z2_L6D4PHI1Z1(
.number_in1(VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1_number),
.read_add1(VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1_read_add),
.innervmstubin(VMS_L5D3PHI1Z2n3_TE_L5D3PHI1Z2_L6D4PHI1Z1),
.number_in2(VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1_number),
.read_add2(VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1_read_add),
.outervmstubin(VMS_L6D4PHI1Z1n1_TE_L5D3PHI1Z2_L6D4PHI1Z1),
.stubpairout(TE_L5D3PHI1Z2_L6D4PHI1Z1_SP_L5D3PHI1Z2_L6D4PHI1Z1),
.valid_data(TE_L5D3PHI1Z2_L6D4PHI1Z1_SP_L5D3PHI1Z2_L6D4PHI1Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI1Z2_L6D4PHI2Z1_phi.txt","TETable_TE_L5D3PHI1Z2_L6D4PHI2Z1_z.txt") TE_L5D3PHI1Z2_L6D4PHI2Z1(
.number_in1(VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1_number),
.read_add1(VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1_read_add),
.innervmstubin(VMS_L5D3PHI1Z2n4_TE_L5D3PHI1Z2_L6D4PHI2Z1),
.number_in2(VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1_number),
.read_add2(VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1_read_add),
.outervmstubin(VMS_L6D4PHI2Z1n1_TE_L5D3PHI1Z2_L6D4PHI2Z1),
.stubpairout(TE_L5D3PHI1Z2_L6D4PHI2Z1_SP_L5D3PHI1Z2_L6D4PHI2Z1),
.valid_data(TE_L5D3PHI1Z2_L6D4PHI2Z1_SP_L5D3PHI1Z2_L6D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI2Z2_L6D4PHI2Z1_phi.txt","TETable_TE_L5D3PHI2Z2_L6D4PHI2Z1_z.txt") TE_L5D3PHI2Z2_L6D4PHI2Z1(
.number_in1(VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1_number),
.read_add1(VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1_read_add),
.innervmstubin(VMS_L5D3PHI2Z2n3_TE_L5D3PHI2Z2_L6D4PHI2Z1),
.number_in2(VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1_number),
.read_add2(VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1_read_add),
.outervmstubin(VMS_L6D4PHI2Z1n2_TE_L5D3PHI2Z2_L6D4PHI2Z1),
.stubpairout(TE_L5D3PHI2Z2_L6D4PHI2Z1_SP_L5D3PHI2Z2_L6D4PHI2Z1),
.valid_data(TE_L5D3PHI2Z2_L6D4PHI2Z1_SP_L5D3PHI2Z2_L6D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI2Z2_L6D4PHI3Z1_phi.txt","TETable_TE_L5D3PHI2Z2_L6D4PHI3Z1_z.txt") TE_L5D3PHI2Z2_L6D4PHI3Z1(
.number_in1(VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1_number),
.read_add1(VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1_read_add),
.innervmstubin(VMS_L5D3PHI2Z2n4_TE_L5D3PHI2Z2_L6D4PHI3Z1),
.number_in2(VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1_number),
.read_add2(VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1_read_add),
.outervmstubin(VMS_L6D4PHI3Z1n1_TE_L5D3PHI2Z2_L6D4PHI3Z1),
.stubpairout(TE_L5D3PHI2Z2_L6D4PHI3Z1_SP_L5D3PHI2Z2_L6D4PHI3Z1),
.valid_data(TE_L5D3PHI2Z2_L6D4PHI3Z1_SP_L5D3PHI2Z2_L6D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI3Z2_L6D4PHI3Z1_phi.txt","TETable_TE_L5D3PHI3Z2_L6D4PHI3Z1_z.txt") TE_L5D3PHI3Z2_L6D4PHI3Z1(
.number_in1(VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1_number),
.read_add1(VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1_read_add),
.innervmstubin(VMS_L5D3PHI3Z2n3_TE_L5D3PHI3Z2_L6D4PHI3Z1),
.number_in2(VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1_number),
.read_add2(VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1_read_add),
.outervmstubin(VMS_L6D4PHI3Z1n2_TE_L5D3PHI3Z2_L6D4PHI3Z1),
.stubpairout(TE_L5D3PHI3Z2_L6D4PHI3Z1_SP_L5D3PHI3Z2_L6D4PHI3Z1),
.valid_data(TE_L5D3PHI3Z2_L6D4PHI3Z1_SP_L5D3PHI3Z2_L6D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D3PHI3Z2_L6D4PHI4Z1_phi.txt","TETable_TE_L5D3PHI3Z2_L6D4PHI4Z1_z.txt") TE_L5D3PHI3Z2_L6D4PHI4Z1(
.number_in1(VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1_number),
.read_add1(VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1_read_add),
.innervmstubin(VMS_L5D3PHI3Z2n4_TE_L5D3PHI3Z2_L6D4PHI4Z1),
.number_in2(VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1_number),
.read_add2(VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1_read_add),
.outervmstubin(VMS_L6D4PHI4Z1n1_TE_L5D3PHI3Z2_L6D4PHI4Z1),
.stubpairout(TE_L5D3PHI3Z2_L6D4PHI4Z1_SP_L5D3PHI3Z2_L6D4PHI4Z1),
.valid_data(TE_L5D3PHI3Z2_L6D4PHI4Z1_SP_L5D3PHI3Z2_L6D4PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI1Z1_L6D4PHI1Z1_phi.txt","TETable_TE_L5D4PHI1Z1_L6D4PHI1Z1_z.txt") TE_L5D4PHI1Z1_L6D4PHI1Z1(
.number_in1(VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1_number),
.read_add1(VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1_read_add),
.outervmstubin(VMS_L6D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI1Z1),
.number_in2(VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1_number),
.read_add2(VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1_read_add),
.innervmstubin(VMS_L5D4PHI1Z1n1_TE_L5D4PHI1Z1_L6D4PHI1Z1),
.stubpairout(TE_L5D4PHI1Z1_L6D4PHI1Z1_SP_L5D4PHI1Z1_L6D4PHI1Z1),
.valid_data(TE_L5D4PHI1Z1_L6D4PHI1Z1_SP_L5D4PHI1Z1_L6D4PHI1Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI1Z1_L6D4PHI2Z1_phi.txt","TETable_TE_L5D4PHI1Z1_L6D4PHI2Z1_z.txt") TE_L5D4PHI1Z1_L6D4PHI2Z1(
.number_in1(VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1_number),
.read_add1(VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1_read_add),
.outervmstubin(VMS_L6D4PHI2Z1n3_TE_L5D4PHI1Z1_L6D4PHI2Z1),
.number_in2(VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1_number),
.read_add2(VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1_read_add),
.innervmstubin(VMS_L5D4PHI1Z1n2_TE_L5D4PHI1Z1_L6D4PHI2Z1),
.stubpairout(TE_L5D4PHI1Z1_L6D4PHI2Z1_SP_L5D4PHI1Z1_L6D4PHI2Z1),
.valid_data(TE_L5D4PHI1Z1_L6D4PHI2Z1_SP_L5D4PHI1Z1_L6D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI2Z1_L6D4PHI2Z1_phi.txt","TETable_TE_L5D4PHI2Z1_L6D4PHI2Z1_z.txt") TE_L5D4PHI2Z1_L6D4PHI2Z1(
.number_in1(VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1_number),
.read_add1(VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1_read_add),
.outervmstubin(VMS_L6D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI2Z1),
.number_in2(VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1_number),
.read_add2(VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1_read_add),
.innervmstubin(VMS_L5D4PHI2Z1n1_TE_L5D4PHI2Z1_L6D4PHI2Z1),
.stubpairout(TE_L5D4PHI2Z1_L6D4PHI2Z1_SP_L5D4PHI2Z1_L6D4PHI2Z1),
.valid_data(TE_L5D4PHI2Z1_L6D4PHI2Z1_SP_L5D4PHI2Z1_L6D4PHI2Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI2Z1_L6D4PHI3Z1_phi.txt","TETable_TE_L5D4PHI2Z1_L6D4PHI3Z1_z.txt") TE_L5D4PHI2Z1_L6D4PHI3Z1(
.number_in1(VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1_number),
.read_add1(VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1_read_add),
.outervmstubin(VMS_L6D4PHI3Z1n3_TE_L5D4PHI2Z1_L6D4PHI3Z1),
.number_in2(VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1_number),
.read_add2(VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1_read_add),
.innervmstubin(VMS_L5D4PHI2Z1n2_TE_L5D4PHI2Z1_L6D4PHI3Z1),
.stubpairout(TE_L5D4PHI2Z1_L6D4PHI3Z1_SP_L5D4PHI2Z1_L6D4PHI3Z1),
.valid_data(TE_L5D4PHI2Z1_L6D4PHI3Z1_SP_L5D4PHI2Z1_L6D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI3Z1_L6D4PHI3Z1_phi.txt","TETable_TE_L5D4PHI3Z1_L6D4PHI3Z1_z.txt") TE_L5D4PHI3Z1_L6D4PHI3Z1(
.number_in1(VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1_number),
.read_add1(VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1_read_add),
.outervmstubin(VMS_L6D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI3Z1),
.number_in2(VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1_number),
.read_add2(VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1_read_add),
.innervmstubin(VMS_L5D4PHI3Z1n1_TE_L5D4PHI3Z1_L6D4PHI3Z1),
.stubpairout(TE_L5D4PHI3Z1_L6D4PHI3Z1_SP_L5D4PHI3Z1_L6D4PHI3Z1),
.valid_data(TE_L5D4PHI3Z1_L6D4PHI3Z1_SP_L5D4PHI3Z1_L6D4PHI3Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI3Z1_L6D4PHI4Z1_phi.txt","TETable_TE_L5D4PHI3Z1_L6D4PHI4Z1_z.txt") TE_L5D4PHI3Z1_L6D4PHI4Z1(
.number_in1(VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_number),
.read_add1(VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_read_add),
.outervmstubin(VMS_L6D4PHI4Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1),
.number_in2(VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_number),
.read_add2(VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1_read_add),
.innervmstubin(VMS_L5D4PHI3Z1n2_TE_L5D4PHI3Z1_L6D4PHI4Z1),
.stubpairout(TE_L5D4PHI3Z1_L6D4PHI4Z1_SP_L5D4PHI3Z1_L6D4PHI4Z1),
.valid_data(TE_L5D4PHI3Z1_L6D4PHI4Z1_SP_L5D4PHI3Z1_L6D4PHI4Z1_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI1Z1_L6D4PHI1Z2_phi.txt","TETable_TE_L5D4PHI1Z1_L6D4PHI1Z2_z.txt") TE_L5D4PHI1Z1_L6D4PHI1Z2(
.number_in1(VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2_number),
.read_add1(VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2_read_add),
.innervmstubin(VMS_L5D4PHI1Z1n3_TE_L5D4PHI1Z1_L6D4PHI1Z2),
.number_in2(VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2_number),
.read_add2(VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2_read_add),
.outervmstubin(VMS_L6D4PHI1Z2n1_TE_L5D4PHI1Z1_L6D4PHI1Z2),
.stubpairout(TE_L5D4PHI1Z1_L6D4PHI1Z2_SP_L5D4PHI1Z1_L6D4PHI1Z2),
.valid_data(TE_L5D4PHI1Z1_L6D4PHI1Z2_SP_L5D4PHI1Z1_L6D4PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI1Z1_L6D4PHI2Z2_phi.txt","TETable_TE_L5D4PHI1Z1_L6D4PHI2Z2_z.txt") TE_L5D4PHI1Z1_L6D4PHI2Z2(
.number_in1(VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2_number),
.read_add1(VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2_read_add),
.innervmstubin(VMS_L5D4PHI1Z1n4_TE_L5D4PHI1Z1_L6D4PHI2Z2),
.number_in2(VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2_number),
.read_add2(VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2_read_add),
.outervmstubin(VMS_L6D4PHI2Z2n1_TE_L5D4PHI1Z1_L6D4PHI2Z2),
.stubpairout(TE_L5D4PHI1Z1_L6D4PHI2Z2_SP_L5D4PHI1Z1_L6D4PHI2Z2),
.valid_data(TE_L5D4PHI1Z1_L6D4PHI2Z2_SP_L5D4PHI1Z1_L6D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI2Z1_L6D4PHI2Z2_phi.txt","TETable_TE_L5D4PHI2Z1_L6D4PHI2Z2_z.txt") TE_L5D4PHI2Z1_L6D4PHI2Z2(
.number_in1(VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2_number),
.read_add1(VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2_read_add),
.innervmstubin(VMS_L5D4PHI2Z1n3_TE_L5D4PHI2Z1_L6D4PHI2Z2),
.number_in2(VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2_number),
.read_add2(VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2_read_add),
.outervmstubin(VMS_L6D4PHI2Z2n2_TE_L5D4PHI2Z1_L6D4PHI2Z2),
.stubpairout(TE_L5D4PHI2Z1_L6D4PHI2Z2_SP_L5D4PHI2Z1_L6D4PHI2Z2),
.valid_data(TE_L5D4PHI2Z1_L6D4PHI2Z2_SP_L5D4PHI2Z1_L6D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI2Z1_L6D4PHI3Z2_phi.txt","TETable_TE_L5D4PHI2Z1_L6D4PHI3Z2_z.txt") TE_L5D4PHI2Z1_L6D4PHI3Z2(
.number_in1(VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2_number),
.read_add1(VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2_read_add),
.innervmstubin(VMS_L5D4PHI2Z1n4_TE_L5D4PHI2Z1_L6D4PHI3Z2),
.number_in2(VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2_number),
.read_add2(VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2_read_add),
.outervmstubin(VMS_L6D4PHI3Z2n1_TE_L5D4PHI2Z1_L6D4PHI3Z2),
.stubpairout(TE_L5D4PHI2Z1_L6D4PHI3Z2_SP_L5D4PHI2Z1_L6D4PHI3Z2),
.valid_data(TE_L5D4PHI2Z1_L6D4PHI3Z2_SP_L5D4PHI2Z1_L6D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI3Z1_L6D4PHI3Z2_phi.txt","TETable_TE_L5D4PHI3Z1_L6D4PHI3Z2_z.txt") TE_L5D4PHI3Z1_L6D4PHI3Z2(
.number_in1(VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2_number),
.read_add1(VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2_read_add),
.innervmstubin(VMS_L5D4PHI3Z1n3_TE_L5D4PHI3Z1_L6D4PHI3Z2),
.number_in2(VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2_number),
.read_add2(VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2_read_add),
.outervmstubin(VMS_L6D4PHI3Z2n2_TE_L5D4PHI3Z1_L6D4PHI3Z2),
.stubpairout(TE_L5D4PHI3Z1_L6D4PHI3Z2_SP_L5D4PHI3Z1_L6D4PHI3Z2),
.valid_data(TE_L5D4PHI3Z1_L6D4PHI3Z2_SP_L5D4PHI3Z1_L6D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI3Z1_L6D4PHI4Z2_phi.txt","TETable_TE_L5D4PHI3Z1_L6D4PHI4Z2_z.txt") TE_L5D4PHI3Z1_L6D4PHI4Z2(
.number_in1(VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2_number),
.read_add1(VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2_read_add),
.innervmstubin(VMS_L5D4PHI3Z1n4_TE_L5D4PHI3Z1_L6D4PHI4Z2),
.number_in2(VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2_number),
.read_add2(VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2_read_add),
.outervmstubin(VMS_L6D4PHI4Z2n1_TE_L5D4PHI3Z1_L6D4PHI4Z2),
.stubpairout(TE_L5D4PHI3Z1_L6D4PHI4Z2_SP_L5D4PHI3Z1_L6D4PHI4Z2),
.valid_data(TE_L5D4PHI3Z1_L6D4PHI4Z2_SP_L5D4PHI3Z1_L6D4PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI1Z2_L6D4PHI1Z2_phi.txt","TETable_TE_L5D4PHI1Z2_L6D4PHI1Z2_z.txt") TE_L5D4PHI1Z2_L6D4PHI1Z2(
.number_in1(VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2_number),
.read_add1(VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2_read_add),
.outervmstubin(VMS_L6D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI1Z2),
.number_in2(VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2_number),
.read_add2(VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2_read_add),
.innervmstubin(VMS_L5D4PHI1Z2n1_TE_L5D4PHI1Z2_L6D4PHI1Z2),
.stubpairout(TE_L5D4PHI1Z2_L6D4PHI1Z2_SP_L5D4PHI1Z2_L6D4PHI1Z2),
.valid_data(TE_L5D4PHI1Z2_L6D4PHI1Z2_SP_L5D4PHI1Z2_L6D4PHI1Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI1Z2_L6D4PHI2Z2_phi.txt","TETable_TE_L5D4PHI1Z2_L6D4PHI2Z2_z.txt") TE_L5D4PHI1Z2_L6D4PHI2Z2(
.number_in1(VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2_number),
.read_add1(VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2_read_add),
.outervmstubin(VMS_L6D4PHI2Z2n3_TE_L5D4PHI1Z2_L6D4PHI2Z2),
.number_in2(VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2_number),
.read_add2(VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2_read_add),
.innervmstubin(VMS_L5D4PHI1Z2n2_TE_L5D4PHI1Z2_L6D4PHI2Z2),
.stubpairout(TE_L5D4PHI1Z2_L6D4PHI2Z2_SP_L5D4PHI1Z2_L6D4PHI2Z2),
.valid_data(TE_L5D4PHI1Z2_L6D4PHI2Z2_SP_L5D4PHI1Z2_L6D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI2Z2_L6D4PHI2Z2_phi.txt","TETable_TE_L5D4PHI2Z2_L6D4PHI2Z2_z.txt") TE_L5D4PHI2Z2_L6D4PHI2Z2(
.number_in1(VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2_number),
.read_add1(VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2_read_add),
.outervmstubin(VMS_L6D4PHI2Z2n4_TE_L5D4PHI2Z2_L6D4PHI2Z2),
.number_in2(VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2_number),
.read_add2(VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2_read_add),
.innervmstubin(VMS_L5D4PHI2Z2n1_TE_L5D4PHI2Z2_L6D4PHI2Z2),
.stubpairout(TE_L5D4PHI2Z2_L6D4PHI2Z2_SP_L5D4PHI2Z2_L6D4PHI2Z2),
.valid_data(TE_L5D4PHI2Z2_L6D4PHI2Z2_SP_L5D4PHI2Z2_L6D4PHI2Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI2Z2_L6D4PHI3Z2_phi.txt","TETable_TE_L5D4PHI2Z2_L6D4PHI3Z2_z.txt") TE_L5D4PHI2Z2_L6D4PHI3Z2(
.number_in1(VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2_number),
.read_add1(VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2_read_add),
.outervmstubin(VMS_L6D4PHI3Z2n3_TE_L5D4PHI2Z2_L6D4PHI3Z2),
.number_in2(VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2_number),
.read_add2(VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2_read_add),
.innervmstubin(VMS_L5D4PHI2Z2n2_TE_L5D4PHI2Z2_L6D4PHI3Z2),
.stubpairout(TE_L5D4PHI2Z2_L6D4PHI3Z2_SP_L5D4PHI2Z2_L6D4PHI3Z2),
.valid_data(TE_L5D4PHI2Z2_L6D4PHI3Z2_SP_L5D4PHI2Z2_L6D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI3Z2_L6D4PHI3Z2_phi.txt","TETable_TE_L5D4PHI3Z2_L6D4PHI3Z2_z.txt") TE_L5D4PHI3Z2_L6D4PHI3Z2(
.number_in1(VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2_number),
.read_add1(VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2_read_add),
.outervmstubin(VMS_L6D4PHI3Z2n4_TE_L5D4PHI3Z2_L6D4PHI3Z2),
.number_in2(VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2_number),
.read_add2(VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2_read_add),
.innervmstubin(VMS_L5D4PHI3Z2n1_TE_L5D4PHI3Z2_L6D4PHI3Z2),
.stubpairout(TE_L5D4PHI3Z2_L6D4PHI3Z2_SP_L5D4PHI3Z2_L6D4PHI3Z2),
.valid_data(TE_L5D4PHI3Z2_L6D4PHI3Z2_SP_L5D4PHI3Z2_L6D4PHI3Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletEngine #("TETable_TE_L5D4PHI3Z2_L6D4PHI4Z2_phi.txt","TETable_TE_L5D4PHI3Z2_L6D4PHI4Z2_z.txt") TE_L5D4PHI3Z2_L6D4PHI4Z2(
.number_in1(VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_number),
.read_add1(VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_read_add),
.outervmstubin(VMS_L6D4PHI4Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2),
.number_in2(VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_number),
.read_add2(VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2_read_add),
.innervmstubin(VMS_L5D4PHI3Z2n2_TE_L5D4PHI3Z2_L6D4PHI4Z2),
.stubpairout(TE_L5D4PHI3Z2_L6D4PHI4Z2_SP_L5D4PHI3Z2_L6D4PHI4Z2),
.valid_data(TE_L5D4PHI3Z2_L6D4PHI4Z2_SP_L5D4PHI3Z2_L6D4PHI4Z2_wr_en),
.start(start3_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator #("InvRTable_TC_L1D3L2D3.dat",`TC_L1L2_krA,`TC_L1L2_krB,1'b1,1'b1) TC_L1D3L2D3(
.number_in1(SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3_number),
.read_add1(SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3_read_add),
.stubpair1in(SP_L1D3PHI1Z1_L2D3PHI1Z1_TC_L1D3L2D3),
.number_in2(SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3_number),
.read_add2(SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3_read_add),
.stubpair2in(SP_L1D3PHI1Z1_L2D3PHI2Z1_TC_L1D3L2D3),
.number_in3(SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3_number),
.read_add3(SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3_read_add),
.stubpair3in(SP_L1D3PHI2Z1_L2D3PHI2Z1_TC_L1D3L2D3),
.number_in4(SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3_number),
.read_add4(SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3_read_add),
.stubpair4in(SP_L1D3PHI2Z1_L2D3PHI3Z1_TC_L1D3L2D3),
.number_in5(SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3_number),
.read_add5(SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3_read_add),
.stubpair5in(SP_L1D3PHI3Z1_L2D3PHI3Z1_TC_L1D3L2D3),
.number_in6(SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3_number),
.read_add6(SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3_read_add),
.stubpair6in(SP_L1D3PHI3Z1_L2D3PHI4Z1_TC_L1D3L2D3),
.number_in7(SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3_number),
.read_add7(SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3_read_add),
.stubpair7in(SP_L1D3PHI1Z1_L2D3PHI1Z2_TC_L1D3L2D3),
.number_in8(SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3_number),
.read_add8(SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3_read_add),
.stubpair8in(SP_L1D3PHI1Z1_L2D3PHI2Z2_TC_L1D3L2D3),
.number_in9(SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3_number),
.read_add9(SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3_read_add),
.stubpair9in(SP_L1D3PHI2Z1_L2D3PHI2Z2_TC_L1D3L2D3),
.number_in10(SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3_number),
.read_add10(SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3_read_add),
.stubpair10in(SP_L1D3PHI2Z1_L2D3PHI3Z2_TC_L1D3L2D3),
.number_in11(SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3_number),
.read_add11(SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3_read_add),
.stubpair11in(SP_L1D3PHI3Z1_L2D3PHI3Z2_TC_L1D3L2D3),
.number_in12(SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3_number),
.read_add12(SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3_read_add),
.stubpair12in(SP_L1D3PHI3Z1_L2D3PHI4Z2_TC_L1D3L2D3),
.number_in13(SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3_number),
.read_add13(SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3_read_add),
.stubpair13in(SP_L1D3PHI1Z2_L2D3PHI1Z2_TC_L1D3L2D3),
.number_in14(SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3_number),
.read_add14(SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3_read_add),
.stubpair14in(SP_L1D3PHI1Z2_L2D3PHI2Z2_TC_L1D3L2D3),
.number_in15(SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3_number),
.read_add15(SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3_read_add),
.stubpair15in(SP_L1D3PHI2Z2_L2D3PHI2Z2_TC_L1D3L2D3),
.number_in16(SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3_number),
.read_add16(SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3_read_add),
.stubpair16in(SP_L1D3PHI2Z2_L2D3PHI3Z2_TC_L1D3L2D3),
.number_in17(SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3_number),
.read_add17(SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3_read_add),
.stubpair17in(SP_L1D3PHI3Z2_L2D3PHI3Z2_TC_L1D3L2D3),
.number_in18(SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3_number),
.read_add18(SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3_read_add),
.stubpair18in(SP_L1D3PHI3Z2_L2D3PHI4Z2_TC_L1D3L2D3),
.read_add_innerall(AS_L1D3n1_TC_L1D3L2D3_read_add),
.innerallstubin(AS_L1D3n1_TC_L1D3L2D3),
.read_add_outerall(AS_L2D3n1_TC_L1D3L2D3_read_add),
.outerallstubin(AS_L2D3n1_TC_L1D3L2D3),
.projoutToPlus_L3(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3),
.projoutToPlus_L4(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4),
.projoutToPlus_L5(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5),
.projoutToPlus_L6(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6),
.projoutToMinus_L3(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3),
.projoutToMinus_L4(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4),
.projoutToMinus_L5(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5),
.projoutToMinus_L6(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6),
.projout_L3D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3),
.projout_L3D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4),
.projout_L4D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3),
.projout_L4D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4),
.projout_L5D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3),
.projout_L5D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4),
.projout_L6D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3),
.projout_L6D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4),
.trackpar(TC_L1D3L2D3_TPAR_L1D3L2D3),
.valid_projoutToPlus_L3(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3_wr_en),
.valid_projoutToPlus_L4(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4_wr_en),
.valid_projoutToPlus_L5(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5_wr_en),
.valid_projoutToPlus_L6(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6_wr_en),
.valid_projoutToMinus_L3(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3_wr_en),
.valid_projoutToMinus_L4(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4_wr_en),
.valid_projoutToMinus_L5(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5_wr_en),
.valid_projoutToMinus_L6(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6_wr_en),
.valid_projout_L3D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3_wr_en),
.valid_projout_L3D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4_wr_en),
.valid_projout_L4D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3_wr_en),
.valid_projout_L4D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4_wr_en),
.valid_projout_L5D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3_wr_en),
.valid_projout_L5D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4_wr_en),
.valid_projout_L6D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3_wr_en),
.valid_projout_L6D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4_wr_en),
.valid_trackpar(TC_L1D3L2D3_TPAR_L1D3L2D3_wr_en),
.done_proj(done_proj4_0),
.start(start4_5),
.done(done4_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator #("InvRTable_TC_L1D3L2D3.dat",`TC_L1L2_krA,`TC_L1L2_krB,1'b1,1'b1)  TC_L1D3L2D4(
.read_add_innerall(AS_L1D3n2_TC_L1D3L2D4_read_add),
.innerallstubin(AS_L1D3n2_TC_L1D3L2D4),
.number_in2(SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4_number),
.read_add2(SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4_read_add),
.stubpair1in(SP_L1D3PHI1Z1_L2D4PHI1Z1_TC_L1D3L2D4),
.number_in3(SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4_number),
.read_add3(SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4_read_add),
.stubpair2in(SP_L1D3PHI1Z1_L2D4PHI2Z1_TC_L1D3L2D4),
.number_in4(SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4_number),
.read_add4(SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4_read_add),
.stubpair3in(SP_L1D3PHI2Z1_L2D4PHI2Z1_TC_L1D3L2D4),
.number_in5(SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4_number),
.read_add5(SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4_read_add),
.stubpair4in(SP_L1D3PHI2Z1_L2D4PHI3Z1_TC_L1D3L2D4),
.number_in6(SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4_number),
.read_add6(SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4_read_add),
.stubpair5in(SP_L1D3PHI3Z1_L2D4PHI3Z1_TC_L1D3L2D4),
.number_in7(SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4_number),
.read_add7(SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4_read_add),
.stubpair6in(SP_L1D3PHI3Z1_L2D4PHI4Z1_TC_L1D3L2D4),
.number_in8(SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4_number),
.read_add8(SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4_read_add),
.stubpair7in(SP_L1D3PHI1Z2_L2D4PHI1Z1_TC_L1D3L2D4),
.number_in9(SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4_number),
.read_add9(SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4_read_add),
.stubpair8in(SP_L1D3PHI1Z2_L2D4PHI2Z1_TC_L1D3L2D4),
.number_in10(SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4_number),
.read_add10(SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4_read_add),
.stubpair9in(SP_L1D3PHI2Z2_L2D4PHI2Z1_TC_L1D3L2D4),
.number_in11(SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4_number),
.read_add11(SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4_read_add),
.stubpair10in(SP_L1D3PHI2Z2_L2D4PHI3Z1_TC_L1D3L2D4),
.number_in12(SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4_number),
.read_add12(SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4_read_add),
.stubpair11in(SP_L1D3PHI3Z2_L2D4PHI3Z1_TC_L1D3L2D4),
.number_in13(SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4_number),
.read_add13(SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4_read_add),
.stubpair12in(SP_L1D3PHI3Z2_L2D4PHI4Z1_TC_L1D3L2D4),
.number_in14(SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4_number),
.read_add14(SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4_read_add),
.stubpair13in(SP_L1D3PHI1Z2_L2D4PHI1Z2_TC_L1D3L2D4),
.number_in15(SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4_number),
.read_add15(SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4_read_add),
.stubpair14in(SP_L1D3PHI1Z2_L2D4PHI2Z2_TC_L1D3L2D4),
.number_in16(SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4_number),
.read_add16(SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4_read_add),
.stubpair15in(SP_L1D3PHI2Z2_L2D4PHI2Z2_TC_L1D3L2D4),
.number_in17(SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4_number),
.read_add17(SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4_read_add),
.stubpair16in(SP_L1D3PHI2Z2_L2D4PHI3Z2_TC_L1D3L2D4),
.number_in18(SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4_number),
.read_add18(SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4_read_add),
.stubpair17in(SP_L1D3PHI3Z2_L2D4PHI3Z2_TC_L1D3L2D4),
.number_in19(SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4_number),
.read_add19(SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4_read_add),
.stubpair18in(SP_L1D3PHI3Z2_L2D4PHI4Z2_TC_L1D3L2D4),
.read_add_outerall(AS_L2D4n1_TC_L1D3L2D4_read_add),
.outerallstubin(AS_L2D4n1_TC_L1D3L2D4),
.projoutToPlus_L3(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3),
.projoutToPlus_L4(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4),
.projoutToPlus_L5(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L5),
.projoutToPlus_L6(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L6),
.projoutToMinus_L3(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3),
.projoutToMinus_L4(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4),
.projoutToMinus_L5(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L5),
.projoutToMinus_L6(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L6),
.projout_L3D3(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D3),
.projout_L3D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4),
.projout_L4D3(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D3),
.projout_L4D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4),
.projout_L5D3(TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D3),
.projout_L5D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D4),
.projout_L6D3(TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D3),
.projout_L6D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D4),
.trackpar(TC_L1D3L2D4_TPAR_L1D3L2D4),
.valid_projoutToPlus_L3(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3_wr_en),
.valid_projoutToPlus_L4(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4_wr_en),
.valid_projoutToPlus_L5(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L5_wr_en),
.valid_projoutToPlus_L6(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L6_wr_en),
.valid_projoutToMinus_L3(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3_wr_en),
.valid_projoutToMinus_L4(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4_wr_en),
.valid_projoutToMinus_L5(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L5_wr_en),
.valid_projoutToMinus_L6(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L6_wr_en),
.valid_projout_L3D3(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D3_wr_en),
.valid_projout_L3D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4_wr_en),
.valid_projout_L4D3(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D3_wr_en),
.valid_projout_L4D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4_wr_en),
.valid_projout_L5D3(TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D3_wr_en),
.valid_projout_L5D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L5D4_wr_en),
.valid_projout_L6D3(TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D3_wr_en),
.valid_projout_L6D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L6D4_wr_en),
.valid_trackpar(TC_L1D3L2D4_TPAR_L1D3L2D4_wr_en),
.start(start4_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator  #("InvRTable_TC_L1D3L2D3.dat",`TC_L1L2_krA,`TC_L1L2_krB,1'b1,1'b1) TC_L1D4L2D4(
.read_add_outerall(AS_L2D4n2_TC_L1D4L2D4_read_add),
.outerallstubin(AS_L2D4n2_TC_L1D4L2D4),
.number_in2(SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4_number),
.read_add2(SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4_read_add),
.stubpair1in(SP_L1D4PHI1Z1_L2D4PHI1Z2_TC_L1D4L2D4),
.number_in3(SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4_number),
.read_add3(SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4_read_add),
.stubpair2in(SP_L1D4PHI1Z1_L2D4PHI2Z2_TC_L1D4L2D4),
.number_in4(SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4_number),
.read_add4(SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4_read_add),
.stubpair3in(SP_L1D4PHI2Z1_L2D4PHI2Z2_TC_L1D4L2D4),
.number_in5(SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4_number),
.read_add5(SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4_read_add),
.stubpair4in(SP_L1D4PHI2Z1_L2D4PHI3Z2_TC_L1D4L2D4),
.number_in6(SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4_number),
.read_add6(SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4_read_add),
.stubpair5in(SP_L1D4PHI3Z1_L2D4PHI3Z2_TC_L1D4L2D4),
.number_in7(SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4_number),
.read_add7(SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4_read_add),
.stubpair6in(SP_L1D4PHI3Z1_L2D4PHI4Z2_TC_L1D4L2D4),
.read_add_innerall(AS_L1D4n1_TC_L1D4L2D4_read_add),
.innerallstubin(AS_L1D4n1_TC_L1D4L2D4),
.projoutToPlus_L3(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3),
.projoutToPlus_L4(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L4),
.projoutToPlus_L5(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L5),
.projoutToPlus_L6(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L6),
.projoutToMinus_L3(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3),
.projoutToMinus_L4(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L4),
.projoutToMinus_L5(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L5),
.projoutToMinus_L6(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L6),
.projout_L3D3(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D3),
.projout_L3D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4),
.projout_L4D3(TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D3),
.projout_L4D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D4),
.projout_L5D3(TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D3),
.projout_L5D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D4),
.projout_L6D3(TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D3),
.projout_L6D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D4),
.trackpar(TC_L1D4L2D4_TPAR_L1D4L2D4),
.valid_projoutToPlus_L3(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3_wr_en),
.valid_projoutToPlus_L4(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L4_wr_en),
.valid_projoutToPlus_L5(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L5_wr_en),
.valid_projoutToPlus_L6(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L6_wr_en),
.valid_projoutToMinus_L3(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3_wr_en),
.valid_projoutToMinus_L4(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L4_wr_en),
.valid_projoutToMinus_L5(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L5_wr_en),
.valid_projoutToMinus_L6(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L6_wr_en),
.valid_projout_L3D3(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D3_wr_en),
.valid_projout_L3D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4_wr_en),
.valid_projout_L4D3(TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D3_wr_en),
.valid_projout_L4D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L4D4_wr_en),
.valid_projout_L5D3(TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D3_wr_en),
.valid_projout_L5D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L5D4_wr_en),
.valid_projout_L6D3(TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D3_wr_en),
.valid_projout_L6D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L6D4_wr_en),
.valid_trackpar(TC_L1D4L2D4_TPAR_L1D4L2D4_wr_en),
.start(start4_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator #("InvRTable_TC_L3D3L4D3.dat",`TC_L3L4_krA,`TC_L3L4_krB,1'b1,1'b0) TC_L3D3L4D3(
.number_in1(SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3_number),
.read_add1(SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3_read_add),
.stubpair1in(SP_L3D3PHI1Z1_L4D3PHI1Z1_TC_L3D3L4D3),
.number_in2(SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3_number),
.read_add2(SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3_read_add),
.stubpair2in(SP_L3D3PHI1Z1_L4D3PHI2Z1_TC_L3D3L4D3),
.number_in3(SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3_number),
.read_add3(SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3_read_add),
.stubpair3in(SP_L3D3PHI2Z1_L4D3PHI2Z1_TC_L3D3L4D3),
.number_in4(SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3_number),
.read_add4(SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3_read_add),
.stubpair4in(SP_L3D3PHI2Z1_L4D3PHI3Z1_TC_L3D3L4D3),
.number_in5(SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3_number),
.read_add5(SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3_read_add),
.stubpair5in(SP_L3D3PHI3Z1_L4D3PHI3Z1_TC_L3D3L4D3),
.number_in6(SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3_number),
.read_add6(SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3_read_add),
.stubpair6in(SP_L3D3PHI3Z1_L4D3PHI4Z1_TC_L3D3L4D3),
.number_in7(SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3_number),
.read_add7(SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3_read_add),
.stubpair7in(SP_L3D3PHI1Z1_L4D3PHI1Z2_TC_L3D3L4D3),
.number_in8(SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3_number),
.read_add8(SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3_read_add),
.stubpair8in(SP_L3D3PHI1Z1_L4D3PHI2Z2_TC_L3D3L4D3),
.number_in9(SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3_number),
.read_add9(SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3_read_add),
.stubpair9in(SP_L3D3PHI2Z1_L4D3PHI2Z2_TC_L3D3L4D3),
.number_in10(SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3_number),
.read_add10(SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3_read_add),
.stubpair10in(SP_L3D3PHI2Z1_L4D3PHI3Z2_TC_L3D3L4D3),
.number_in11(SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3_number),
.read_add11(SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3_read_add),
.stubpair11in(SP_L3D3PHI3Z1_L4D3PHI3Z2_TC_L3D3L4D3),
.number_in12(SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3_number),
.read_add12(SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3_read_add),
.stubpair12in(SP_L3D3PHI3Z1_L4D3PHI4Z2_TC_L3D3L4D3),
.number_in13(SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3_number),
.read_add13(SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3_read_add),
.stubpair13in(SP_L3D3PHI1Z2_L4D3PHI1Z2_TC_L3D3L4D3),
.number_in14(SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3_number),
.read_add14(SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3_read_add),
.stubpair14in(SP_L3D3PHI1Z2_L4D3PHI2Z2_TC_L3D3L4D3),
.number_in15(SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3_number),
.read_add15(SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3_read_add),
.stubpair15in(SP_L3D3PHI2Z2_L4D3PHI2Z2_TC_L3D3L4D3),
.number_in16(SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3_number),
.read_add16(SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3_read_add),
.stubpair16in(SP_L3D3PHI2Z2_L4D3PHI3Z2_TC_L3D3L4D3),
.number_in17(SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3_number),
.read_add17(SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3_read_add),
.stubpair17in(SP_L3D3PHI3Z2_L4D3PHI3Z2_TC_L3D3L4D3),
.number_in18(SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3_number),
.read_add18(SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3_read_add),
.stubpair18in(SP_L3D3PHI3Z2_L4D3PHI4Z2_TC_L3D3L4D3),
.read_add_innerall(AS_L3D3n1_TC_L3D3L4D3_read_add),
.innerallstubin(AS_L3D3n1_TC_L3D3L4D3),
.read_add_outerall(AS_L4D3n1_TC_L3D3L4D3_read_add),
.outerallstubin(AS_L4D3n1_TC_L3D3L4D3),
.projoutToPlus_L1(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1),
.projoutToPlus_L2(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2),
.projoutToPlus_L5(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5),
.projoutToPlus_L6(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6),
.projoutToMinus_L1(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1),
.projoutToMinus_L2(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2),
.projoutToMinus_L5(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5),
.projoutToMinus_L6(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6),
.projout_L1D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3),
.projout_L1D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D4),
.projout_L2D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3),
.projout_L2D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D4),
.projout_L5D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3),
.projout_L5D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4),
.projout_L6D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3),
.projout_L6D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4),
.trackpar(TC_L3D3L4D3_TPAR_L3D3L4D3),
.valid_projoutToPlus_L1(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1_wr_en),
.valid_projoutToPlus_L2(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2_wr_en),
.valid_projoutToPlus_L5(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5_wr_en),
.valid_projoutToPlus_L6(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6_wr_en),
.valid_projoutToMinus_L1(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1_wr_en),
.valid_projoutToMinus_L2(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2_wr_en),
.valid_projoutToMinus_L5(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5_wr_en),
.valid_projoutToMinus_L6(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6_wr_en),
.valid_projout_L1D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3_wr_en),
.valid_projout_L1D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D4_wr_en),
.valid_projout_L2D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3_wr_en),
.valid_projout_L2D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D4_wr_en),
.valid_projout_L5D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3_wr_en),
.valid_projout_L5D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4_wr_en),
.valid_projout_L6D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3_wr_en),
.valid_projout_L6D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4_wr_en),
.valid_trackpar(TC_L3D3L4D3_TPAR_L3D3L4D3_wr_en),
.start(start4_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator #("InvRTable_TC_L3D3L4D3.dat",`TC_L3L4_krA,`TC_L3L4_krB,1'b1,1'b0) TC_L3D3L4D4(
.read_add_innerall(AS_L3D3n2_TC_L3D3L4D4_read_add),
.innerallstubin(AS_L3D3n2_TC_L3D3L4D4),
.number_in2(SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4_number),
.read_add2(SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4_read_add),
.stubpair1in(SP_L3D3PHI1Z2_L4D4PHI1Z1_TC_L3D3L4D4),
.number_in3(SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4_number),
.read_add3(SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4_read_add),
.stubpair2in(SP_L3D3PHI1Z2_L4D4PHI2Z1_TC_L3D3L4D4),
.number_in4(SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4_number),
.read_add4(SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4_read_add),
.stubpair3in(SP_L3D3PHI2Z2_L4D4PHI2Z1_TC_L3D3L4D4),
.number_in5(SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4_number),
.read_add5(SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4_read_add),
.stubpair4in(SP_L3D3PHI2Z2_L4D4PHI3Z1_TC_L3D3L4D4),
.number_in6(SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4_number),
.read_add6(SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4_read_add),
.stubpair5in(SP_L3D3PHI3Z2_L4D4PHI3Z1_TC_L3D3L4D4),
.number_in7(SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4_number),
.read_add7(SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4_read_add),
.stubpair6in(SP_L3D3PHI3Z2_L4D4PHI4Z1_TC_L3D3L4D4),
.read_add_outerall(AS_L4D4n1_TC_L3D3L4D4_read_add),
.outerallstubin(AS_L4D4n1_TC_L3D3L4D4),
.projoutToPlus_L1(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1),
.projoutToPlus_L2(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2),
.projoutToPlus_L5(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5),
.projoutToPlus_L6(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6),
.projoutToMinus_L1(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1),
.projoutToMinus_L2(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2),
.projoutToMinus_L5(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5),
.projoutToMinus_L6(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6),
.projout_L1D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3),
.projout_L1D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D4),
.projout_L2D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3),
.projout_L2D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D4),
.projout_L5D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D3),
.projout_L5D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4),
.projout_L6D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D3),
.projout_L6D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4),
.trackpar(TC_L3D3L4D4_TPAR_L3D3L4D4),
.valid_projoutToPlus_L1(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1_wr_en),
.valid_projoutToPlus_L2(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2_wr_en),
.valid_projoutToPlus_L5(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5_wr_en),
.valid_projoutToPlus_L6(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6_wr_en),
.valid_projoutToMinus_L1(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1_wr_en),
.valid_projoutToMinus_L2(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2_wr_en),
.valid_projoutToMinus_L5(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5_wr_en),
.valid_projoutToMinus_L6(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6_wr_en),
.valid_projout_L1D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3_wr_en),
.valid_projout_L1D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D4_wr_en),
.valid_projout_L2D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3_wr_en),
.valid_projout_L2D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D4_wr_en),
.valid_projout_L5D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D3_wr_en),
.valid_projout_L5D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4_wr_en),
.valid_projout_L6D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D3_wr_en),
.valid_projout_L6D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4_wr_en),
.valid_trackpar(TC_L3D3L4D4_TPAR_L3D3L4D4_wr_en),
.start(start4_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator #("InvRTable_TC_L3D3L4D3.dat",`TC_L3L4_krA,`TC_L3L4_krB,1'b1,1'b0) TC_L3D4L4D4(
.read_add_outerall(AS_L4D4n2_TC_L3D4L4D4_read_add),
.outerallstubin(AS_L4D4n2_TC_L3D4L4D4),
.number_in2(SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4_number),
.read_add2(SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4_read_add),
.stubpair1in(SP_L3D4PHI1Z1_L4D4PHI1Z1_TC_L3D4L4D4),
.number_in3(SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4_number),
.read_add3(SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4_read_add),
.stubpair2in(SP_L3D4PHI1Z1_L4D4PHI2Z1_TC_L3D4L4D4),
.number_in4(SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4_number),
.read_add4(SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4_read_add),
.stubpair3in(SP_L3D4PHI2Z1_L4D4PHI2Z1_TC_L3D4L4D4),
.number_in5(SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4_number),
.read_add5(SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4_read_add),
.stubpair4in(SP_L3D4PHI2Z1_L4D4PHI3Z1_TC_L3D4L4D4),
.number_in6(SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4_number),
.read_add6(SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4_read_add),
.stubpair5in(SP_L3D4PHI3Z1_L4D4PHI3Z1_TC_L3D4L4D4),
.number_in7(SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4_number),
.read_add7(SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4_read_add),
.stubpair6in(SP_L3D4PHI3Z1_L4D4PHI4Z1_TC_L3D4L4D4),
.number_in8(SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4_number),
.read_add8(SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4_read_add),
.stubpair7in(SP_L3D4PHI1Z1_L4D4PHI1Z2_TC_L3D4L4D4),
.number_in9(SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4_number),
.read_add9(SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4_read_add),
.stubpair8in(SP_L3D4PHI1Z1_L4D4PHI2Z2_TC_L3D4L4D4),
.number_in10(SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4_number),
.read_add10(SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4_read_add),
.stubpair9in(SP_L3D4PHI2Z1_L4D4PHI2Z2_TC_L3D4L4D4),
.number_in11(SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4_number),
.read_add11(SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4_read_add),
.stubpair10in(SP_L3D4PHI2Z1_L4D4PHI3Z2_TC_L3D4L4D4),
.number_in12(SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4_number),
.read_add12(SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4_read_add),
.stubpair11in(SP_L3D4PHI3Z1_L4D4PHI3Z2_TC_L3D4L4D4),
.number_in13(SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4_number),
.read_add13(SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4_read_add),
.stubpair12in(SP_L3D4PHI3Z1_L4D4PHI4Z2_TC_L3D4L4D4),
.number_in14(SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4_number),
.read_add14(SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4_read_add),
.stubpair13in(SP_L3D4PHI1Z2_L4D4PHI1Z2_TC_L3D4L4D4),
.number_in15(SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4_number),
.read_add15(SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4_read_add),
.stubpair14in(SP_L3D4PHI1Z2_L4D4PHI2Z2_TC_L3D4L4D4),
.number_in16(SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4_number),
.read_add16(SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4_read_add),
.stubpair15in(SP_L3D4PHI2Z2_L4D4PHI2Z2_TC_L3D4L4D4),
.number_in17(SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4_number),
.read_add17(SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4_read_add),
.stubpair16in(SP_L3D4PHI2Z2_L4D4PHI3Z2_TC_L3D4L4D4),
.number_in18(SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4_number),
.read_add18(SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4_read_add),
.stubpair17in(SP_L3D4PHI3Z2_L4D4PHI3Z2_TC_L3D4L4D4),
.number_in19(SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4_number),
.read_add19(SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4_read_add),
.stubpair18in(SP_L3D4PHI3Z2_L4D4PHI4Z2_TC_L3D4L4D4),
.read_add_innerall(AS_L3D4n1_TC_L3D4L4D4_read_add),
.innerallstubin(AS_L3D4n1_TC_L3D4L4D4),
.projoutToPlus_L1(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1),
.projoutToPlus_L2(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2),
.projoutToPlus_L5(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5),
.projoutToPlus_L6(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6),
.projoutToMinus_L1(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1),
.projoutToMinus_L2(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2),
.projoutToMinus_L5(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5),
.projoutToMinus_L6(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6),
.projout_L1D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3),
.projout_L1D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D4),
.projout_L2D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3),
.projout_L2D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4),
.projout_L5D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D3),
.projout_L5D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4),
.projout_L6D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D3),
.projout_L6D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4),
.trackpar(TC_L3D4L4D4_TPAR_L3D4L4D4),
.valid_projoutToPlus_L1(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1_wr_en),
.valid_projoutToPlus_L2(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2_wr_en),
.valid_projoutToPlus_L5(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5_wr_en),
.valid_projoutToPlus_L6(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6_wr_en),
.valid_projoutToMinus_L1(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1_wr_en),
.valid_projoutToMinus_L2(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2_wr_en),
.valid_projoutToMinus_L5(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5_wr_en),
.valid_projoutToMinus_L6(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6_wr_en),
.valid_projout_L1D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3_wr_en),
.valid_projout_L1D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D4_wr_en),
.valid_projout_L2D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3_wr_en),
.valid_projout_L2D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4_wr_en),
.valid_projout_L5D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D3_wr_en),
.valid_projout_L5D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4_wr_en),
.valid_projout_L6D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D3_wr_en),
.valid_projout_L6D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4_wr_en),
.valid_trackpar(TC_L3D4L4D4_TPAR_L3D4L4D4_wr_en),
.start(start4_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator #("InvRTable_TC_L5D3L6D3.dat",`TC_L5L6_krA,`TC_L5L6_krB,1'b0,1'b0) TC_L5D3L6D3(
.number_in1(SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3_number),
.read_add1(SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3_read_add),
.stubpair1in(SP_L5D3PHI1Z1_L6D3PHI1Z1_TC_L5D3L6D3),
.number_in2(SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3_number),
.read_add2(SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3_read_add),
.stubpair2in(SP_L5D3PHI1Z1_L6D3PHI2Z1_TC_L5D3L6D3),
.number_in3(SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3_number),
.read_add3(SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3_read_add),
.stubpair3in(SP_L5D3PHI2Z1_L6D3PHI2Z1_TC_L5D3L6D3),
.number_in4(SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3_number),
.read_add4(SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3_read_add),
.stubpair4in(SP_L5D3PHI2Z1_L6D3PHI3Z1_TC_L5D3L6D3),
.number_in5(SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3_number),
.read_add5(SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3_read_add),
.stubpair5in(SP_L5D3PHI3Z1_L6D3PHI3Z1_TC_L5D3L6D3),
.number_in6(SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3_number),
.read_add6(SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3_read_add),
.stubpair6in(SP_L5D3PHI3Z1_L6D3PHI4Z1_TC_L5D3L6D3),
.number_in7(SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3_number),
.read_add7(SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3_read_add),
.stubpair7in(SP_L5D3PHI1Z1_L6D3PHI1Z2_TC_L5D3L6D3),
.number_in8(SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3_number),
.read_add8(SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3_read_add),
.stubpair8in(SP_L5D3PHI1Z1_L6D3PHI2Z2_TC_L5D3L6D3),
.number_in9(SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3_number),
.read_add9(SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3_read_add),
.stubpair9in(SP_L5D3PHI2Z1_L6D3PHI2Z2_TC_L5D3L6D3),
.number_in10(SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3_number),
.read_add10(SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3_read_add),
.stubpair10in(SP_L5D3PHI2Z1_L6D3PHI3Z2_TC_L5D3L6D3),
.number_in11(SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3_number),
.read_add11(SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3_read_add),
.stubpair11in(SP_L5D3PHI3Z1_L6D3PHI3Z2_TC_L5D3L6D3),
.number_in12(SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3_number),
.read_add12(SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3_read_add),
.stubpair12in(SP_L5D3PHI3Z1_L6D3PHI4Z2_TC_L5D3L6D3),
.number_in13(SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3_number),
.read_add13(SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3_read_add),
.stubpair13in(SP_L5D3PHI1Z2_L6D3PHI1Z2_TC_L5D3L6D3),
.number_in14(SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3_number),
.read_add14(SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3_read_add),
.stubpair14in(SP_L5D3PHI1Z2_L6D3PHI2Z2_TC_L5D3L6D3),
.number_in15(SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3_number),
.read_add15(SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3_read_add),
.stubpair15in(SP_L5D3PHI2Z2_L6D3PHI2Z2_TC_L5D3L6D3),
.number_in16(SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3_number),
.read_add16(SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3_read_add),
.stubpair16in(SP_L5D3PHI2Z2_L6D3PHI3Z2_TC_L5D3L6D3),
.number_in17(SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3_number),
.read_add17(SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3_read_add),
.stubpair17in(SP_L5D3PHI3Z2_L6D3PHI3Z2_TC_L5D3L6D3),
.number_in18(SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3_number),
.read_add18(SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3_read_add),
.stubpair18in(SP_L5D3PHI3Z2_L6D3PHI4Z2_TC_L5D3L6D3),
.read_add_innerall(AS_L5D3n1_TC_L5D3L6D3_read_add),
.innerallstubin(AS_L5D3n1_TC_L5D3L6D3),
.read_add_outerall(AS_L6D3n1_TC_L5D3L6D3_read_add),
.outerallstubin(AS_L6D3n1_TC_L5D3L6D3),
.projoutToPlus_L1(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1),
.projoutToPlus_L2(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2),
.projoutToPlus_L3(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3),
.projoutToPlus_L4(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4),
.projoutToMinus_L1(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1),
.projoutToMinus_L2(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2),
.projoutToMinus_L3(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3),
.projoutToMinus_L4(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4),
.projout_L1D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3),
.projout_L1D4(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D4),
.projout_L2D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3),
.projout_L2D4(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D4),
.projout_L3D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3),
.projout_L3D4(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D4),
.projout_L4D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3),
.projout_L4D4(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D4),
.trackpar(TC_L5D3L6D3_TPAR_L5D3L6D3),
.valid_projoutToPlus_L1(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1_wr_en),
.valid_projoutToPlus_L2(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2_wr_en),
.valid_projoutToPlus_L3(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3_wr_en),
.valid_projoutToPlus_L4(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4_wr_en),
.valid_projoutToMinus_L1(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1_wr_en),
.valid_projoutToMinus_L2(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2_wr_en),
.valid_projoutToMinus_L3(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3_wr_en),
.valid_projoutToMinus_L4(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4_wr_en),
.valid_projout_L1D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3_wr_en),
.valid_projout_L1D4(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D4_wr_en),
.valid_projout_L2D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3_wr_en),
.valid_projout_L2D4(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D4_wr_en),
.valid_projout_L3D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3_wr_en),
.valid_projout_L3D4(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D4_wr_en),
.valid_projout_L4D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3_wr_en),
.valid_projout_L4D4(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D4_wr_en),
.valid_trackpar(TC_L5D3L6D3_TPAR_L5D3L6D3_wr_en),
.start(start4_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator #("InvRTable_TC_L5D3L6D3.dat",`TC_L5L6_krA,`TC_L5L6_krB,1'b0,1'b0) TC_L5D3L6D4(
.read_add_innerall(AS_L5D3n2_TC_L5D3L6D4_read_add),
.innerallstubin(AS_L5D3n2_TC_L5D3L6D4),
.number_in2(SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4_number),
.read_add2(SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4_read_add),
.stubpair1in(SP_L5D3PHI1Z2_L6D4PHI1Z1_TC_L5D3L6D4),
.number_in3(SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4_number),
.read_add3(SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4_read_add),
.stubpair2in(SP_L5D3PHI1Z2_L6D4PHI2Z1_TC_L5D3L6D4),
.number_in4(SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4_number),
.read_add4(SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4_read_add),
.stubpair3in(SP_L5D3PHI2Z2_L6D4PHI2Z1_TC_L5D3L6D4),
.number_in5(SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4_number),
.read_add5(SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4_read_add),
.stubpair4in(SP_L5D3PHI2Z2_L6D4PHI3Z1_TC_L5D3L6D4),
.number_in6(SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4_number),
.read_add6(SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4_read_add),
.stubpair5in(SP_L5D3PHI3Z2_L6D4PHI3Z1_TC_L5D3L6D4),
.number_in7(SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4_number),
.read_add7(SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4_read_add),
.stubpair6in(SP_L5D3PHI3Z2_L6D4PHI4Z1_TC_L5D3L6D4),
.read_add_outerall(AS_L6D4n1_TC_L5D3L6D4_read_add),
.outerallstubin(AS_L6D4n1_TC_L5D3L6D4),
.projoutToPlus_L1(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1),
.projoutToPlus_L2(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2),
.projoutToPlus_L3(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3),
.projoutToPlus_L4(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4),
.projoutToMinus_L1(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1),
.projoutToMinus_L2(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2),
.projoutToMinus_L3(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3),
.projoutToMinus_L4(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4),
.projout_L1D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3),
.projout_L1D4(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D4),
.projout_L2D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3),
.projout_L2D4(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D4),
.projout_L3D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3),
.projout_L3D4(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D4),
.projout_L4D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3),
.projout_L4D4(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D4),
.trackpar(TC_L5D3L6D4_TPAR_L5D3L6D4),
.valid_projoutToPlus_L1(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1_wr_en),
.valid_projoutToPlus_L2(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2_wr_en),
.valid_projoutToPlus_L3(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3_wr_en),
.valid_projoutToPlus_L4(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4_wr_en),
.valid_projoutToMinus_L1(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1_wr_en),
.valid_projoutToMinus_L2(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2_wr_en),
.valid_projoutToMinus_L3(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3_wr_en),
.valid_projoutToMinus_L4(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4_wr_en),
.valid_projout_L1D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3_wr_en),
.valid_projout_L1D4(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D4_wr_en),
.valid_projout_L2D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3_wr_en),
.valid_projout_L2D4(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D4_wr_en),
.valid_projout_L3D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3_wr_en),
.valid_projout_L3D4(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D4_wr_en),
.valid_projout_L4D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3_wr_en),
.valid_projout_L4D4(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D4_wr_en),
.valid_trackpar(TC_L5D3L6D4_TPAR_L5D3L6D4_wr_en),
.start(start4_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


TrackletCalculator #("InvRTable_TC_L5D3L6D3.dat",`TC_L5L6_krA,`TC_L5L6_krB,1'b0,1'b0) TC_L5D4L6D4(
.read_add_outerall(AS_L6D4n2_TC_L5D4L6D4_read_add),
.outerallstubin(AS_L6D4n2_TC_L5D4L6D4),
.number_in2(SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4_number),
.read_add2(SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4_read_add),
.stubpair1in(SP_L5D4PHI1Z1_L6D4PHI1Z1_TC_L5D4L6D4),
.number_in3(SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4_number),
.read_add3(SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4_read_add),
.stubpair2in(SP_L5D4PHI1Z1_L6D4PHI2Z1_TC_L5D4L6D4),
.number_in4(SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4_number),
.read_add4(SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4_read_add),
.stubpair3in(SP_L5D4PHI2Z1_L6D4PHI2Z1_TC_L5D4L6D4),
.number_in5(SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4_number),
.read_add5(SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4_read_add),
.stubpair4in(SP_L5D4PHI2Z1_L6D4PHI3Z1_TC_L5D4L6D4),
.number_in6(SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4_number),
.read_add6(SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4_read_add),
.stubpair5in(SP_L5D4PHI3Z1_L6D4PHI3Z1_TC_L5D4L6D4),
.number_in7(SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4_number),
.read_add7(SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4_read_add),
.stubpair6in(SP_L5D4PHI3Z1_L6D4PHI4Z1_TC_L5D4L6D4),
.number_in8(SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4_number),
.read_add8(SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4_read_add),
.stubpair7in(SP_L5D4PHI1Z1_L6D4PHI1Z2_TC_L5D4L6D4),
.number_in9(SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4_number),
.read_add9(SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4_read_add),
.stubpair8in(SP_L5D4PHI1Z1_L6D4PHI2Z2_TC_L5D4L6D4),
.number_in10(SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4_number),
.read_add10(SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4_read_add),
.stubpair9in(SP_L5D4PHI2Z1_L6D4PHI2Z2_TC_L5D4L6D4),
.number_in11(SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4_number),
.read_add11(SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4_read_add),
.stubpair10in(SP_L5D4PHI2Z1_L6D4PHI3Z2_TC_L5D4L6D4),
.number_in12(SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4_number),
.read_add12(SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4_read_add),
.stubpair11in(SP_L5D4PHI3Z1_L6D4PHI3Z2_TC_L5D4L6D4),
.number_in13(SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4_number),
.read_add13(SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4_read_add),
.stubpair12in(SP_L5D4PHI3Z1_L6D4PHI4Z2_TC_L5D4L6D4),
.number_in14(SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4_number),
.read_add14(SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4_read_add),
.stubpair13in(SP_L5D4PHI1Z2_L6D4PHI1Z2_TC_L5D4L6D4),
.number_in15(SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4_number),
.read_add15(SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4_read_add),
.stubpair14in(SP_L5D4PHI1Z2_L6D4PHI2Z2_TC_L5D4L6D4),
.number_in16(SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4_number),
.read_add16(SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4_read_add),
.stubpair15in(SP_L5D4PHI2Z2_L6D4PHI2Z2_TC_L5D4L6D4),
.number_in17(SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4_number),
.read_add17(SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4_read_add),
.stubpair16in(SP_L5D4PHI2Z2_L6D4PHI3Z2_TC_L5D4L6D4),
.number_in18(SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4_number),
.read_add18(SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4_read_add),
.stubpair17in(SP_L5D4PHI3Z2_L6D4PHI3Z2_TC_L5D4L6D4),
.number_in19(SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4_number),
.read_add19(SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4_read_add),
.stubpair18in(SP_L5D4PHI3Z2_L6D4PHI4Z2_TC_L5D4L6D4),
.read_add_innerall(AS_L5D4n1_TC_L5D4L6D4_read_add),
.innerallstubin(AS_L5D4n1_TC_L5D4L6D4),
.projoutToPlus_L1(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1),
.projoutToPlus_L2(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2),
.projoutToPlus_L3(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3),
.projoutToPlus_L4(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4),
.projoutToMinus_L1(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1),
.projoutToMinus_L2(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2),
.projoutToMinus_L3(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3),
.projoutToMinus_L4(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4),
.projout_L1D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3),
.projout_L1D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D4),
.projout_L2D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3),
.projout_L2D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D4),
.projout_L3D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3),
.projout_L3D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4),
.projout_L4D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3),
.projout_L4D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4),
.trackpar(TC_L5D4L6D4_TPAR_L5D4L6D4),
.valid_projoutToPlus_L1(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1_wr_en),
.valid_projoutToPlus_L2(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2_wr_en),
.valid_projoutToPlus_L3(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3_wr_en),
.valid_projoutToPlus_L4(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4_wr_en),
.valid_projoutToMinus_L1(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1_wr_en),
.valid_projoutToMinus_L2(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2_wr_en),
.valid_projoutToMinus_L3(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3_wr_en),
.valid_projoutToMinus_L4(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4_wr_en),
.valid_projout_L1D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3_wr_en),
.valid_projout_L1D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D4_wr_en),
.valid_projout_L2D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3_wr_en),
.valid_projout_L2D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D4_wr_en),
.valid_projout_L3D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3_wr_en),
.valid_projout_L3D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4_wr_en),
.valid_projout_L4D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3_wr_en),
.valid_projout_L4D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4_wr_en),
.valid_trackpar(TC_L5D4L6D4_TPAR_L5D4L6D4_wr_en),
.start(start4_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionTransceiver  PT_L1L2_Plus(
.number_in1(TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus_number),
.read_add1(TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus_read_add),
.projin_1(TPROJ_ToPlus_L1D3L2D3_L3_PT_L1L2_Plus),
.number_in2(TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus_number),
.read_add2(TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus_read_add),
.projin_2(TPROJ_ToPlus_L1D3L2D3_L4_PT_L1L2_Plus),
.number_in3(TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus_number),
.read_add3(TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus_read_add),
.projin_3(TPROJ_ToPlus_L1D3L2D3_L5_PT_L1L2_Plus),
.number_in4(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus_number),
.read_add4(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus_read_add),
.projin_4(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L2_Plus),
.number_in5(TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus_number),
.read_add5(TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus_read_add),
.projin_5(TPROJ_ToPlus_L1D3L2D4_L3_PT_L1L2_Plus),
.number_in6(TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus_number),
.read_add6(TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus_read_add),
.projin_6(TPROJ_ToPlus_L1D3L2D4_L4_PT_L1L2_Plus),
.number_in7(TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus_number),
.read_add7(TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus_read_add),
.projin_7(TPROJ_ToPlus_L1D3L2D4_L5_PT_L1L2_Plus),
.number_in8(TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus_number),
.read_add8(TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus_read_add),
.projin_8(TPROJ_ToPlus_L1D3L2D4_L6_PT_L1L2_Plus),
.number_in9(TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus_number),
.read_add9(TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus_read_add),
.projin_9(TPROJ_ToPlus_L1D4L2D4_L3_PT_L1L2_Plus),
.number_in10(TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus_number),
.read_add10(TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus_read_add),
.projin_10(TPROJ_ToPlus_L1D4L2D4_L4_PT_L1L2_Plus),
.number_in11(TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus_number),
.read_add11(TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus_read_add),
.projin_11(TPROJ_ToPlus_L1D4L2D4_L5_PT_L1L2_Plus),
.number_in12(TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus_number),
.read_add12(TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus_read_add),
.projin_12(TPROJ_ToPlus_L1D4L2D4_L6_PT_L1L2_Plus),
.valid_incomming_proj_data_stream(PT_L1L2_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L1L2_Plus_From_DataStream),
.projout_1(PT_L1L2_Plus_TPROJ_FromPlus_L3D3_L1L2),
.projout_2(PT_L1L2_Plus_TPROJ_FromPlus_L3D4_L1L2),
.projout_3(PT_L1L2_Plus_TPROJ_FromPlus_L4D3_L1L2),
.projout_4(PT_L1L2_Plus_TPROJ_FromPlus_L4D4_L1L2),
.projout_5(PT_L1L2_Plus_TPROJ_FromPlus_L5D3_L1L2),
.projout_6(PT_L1L2_Plus_TPROJ_FromPlus_L5D4_L1L2),
.projout_7(PT_L1L2_Plus_TPROJ_FromPlus_L6D3_L1L2),
.projout_8(PT_L1L2_Plus_TPROJ_FromPlus_L6D4_L1L2),
.valid_1(PT_L1L2_Plus_TPROJ_FromPlus_L3D3_L1L2_wr_en),
.valid_2(PT_L1L2_Plus_TPROJ_FromPlus_L3D4_L1L2_wr_en),
.valid_3(PT_L1L2_Plus_TPROJ_FromPlus_L4D3_L1L2_wr_en),
.valid_4(PT_L1L2_Plus_TPROJ_FromPlus_L4D4_L1L2_wr_en),
.valid_5(PT_L1L2_Plus_TPROJ_FromPlus_L5D3_L1L2_wr_en),
.valid_6(PT_L1L2_Plus_TPROJ_FromPlus_L5D4_L1L2_wr_en),
.valid_7(PT_L1L2_Plus_TPROJ_FromPlus_L6D3_L1L2_wr_en),
.valid_8(PT_L1L2_Plus_TPROJ_FromPlus_L6D4_L1L2_wr_en),
.valid_proj_data_stream(PT_L1L2_Plus_To_DataStream_en),
.proj_data_stream(PT_L1L2_Plus_To_DataStream),
.start(start5_5),
.done(done5_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionTransceiver  PT_L3L4_Plus(
.number_in1(TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus_number),
.read_add1(TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus_read_add),
.projin_1(TPROJ_ToPlus_L3D3L4D3_L1_PT_L3L4_Plus),
.number_in2(TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus_number),
.read_add2(TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus_read_add),
.projin_2(TPROJ_ToPlus_L3D3L4D3_L2_PT_L3L4_Plus),
.number_in3(TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus_number),
.read_add3(TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus_read_add),
.projin_3(TPROJ_ToPlus_L3D3L4D3_L5_PT_L3L4_Plus),
.number_in4(TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus_number),
.read_add4(TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus_read_add),
.projin_4(TPROJ_ToPlus_L3D3L4D3_L6_PT_L3L4_Plus),
.number_in5(TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus_number),
.read_add5(TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus_read_add),
.projin_5(TPROJ_ToPlus_L3D3L4D4_L1_PT_L3L4_Plus),
.number_in6(TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus_number),
.read_add6(TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus_read_add),
.projin_6(TPROJ_ToPlus_L3D3L4D4_L2_PT_L3L4_Plus),
.number_in7(TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus_number),
.read_add7(TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus_read_add),
.projin_7(TPROJ_ToPlus_L3D3L4D4_L5_PT_L3L4_Plus),
.number_in8(TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus_number),
.read_add8(TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus_read_add),
.projin_8(TPROJ_ToPlus_L3D3L4D4_L6_PT_L3L4_Plus),
.number_in9(TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus_number),
.read_add9(TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus_read_add),
.projin_9(TPROJ_ToPlus_L3D4L4D4_L1_PT_L3L4_Plus),
.number_in10(TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus_number),
.read_add10(TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus_read_add),
.projin_10(TPROJ_ToPlus_L3D4L4D4_L2_PT_L3L4_Plus),
.number_in11(TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus_number),
.read_add11(TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus_read_add),
.projin_11(TPROJ_ToPlus_L3D4L4D4_L5_PT_L3L4_Plus),
.number_in12(TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus_number),
.read_add12(TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus_read_add),
.projin_12(TPROJ_ToPlus_L3D4L4D4_L6_PT_L3L4_Plus),
.valid_incomming_proj_data_stream(PT_L3L4_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L3L4_Plus_From_DataStream),
.projout_1(PT_L3L4_Plus_TPROJ_FromPlus_L1D3_L3L4),
.projout_2(PT_L3L4_Plus_TPROJ_FromPlus_L1D4_L3L4),
.projout_3(PT_L3L4_Plus_TPROJ_FromPlus_L2D3_L3L4),
.projout_4(PT_L3L4_Plus_TPROJ_FromPlus_L2D4_L3L4),
.projout_5(PT_L3L4_Plus_TPROJ_FromPlus_L5D3_L3L4),
.projout_6(PT_L3L4_Plus_TPROJ_FromPlus_L5D4_L3L4),
.projout_7(PT_L3L4_Plus_TPROJ_FromPlus_L6D3_L3L4),
.projout_8(PT_L3L4_Plus_TPROJ_FromPlus_L6D4_L3L4),
.valid_1(PT_L3L4_Plus_TPROJ_FromPlus_L1D3_L3L4_wr_en),
.valid_2(PT_L3L4_Plus_TPROJ_FromPlus_L1D4_L3L4_wr_en),
.valid_3(PT_L3L4_Plus_TPROJ_FromPlus_L2D3_L3L4_wr_en),
.valid_4(PT_L3L4_Plus_TPROJ_FromPlus_L2D4_L3L4_wr_en),
.valid_5(PT_L3L4_Plus_TPROJ_FromPlus_L5D3_L3L4_wr_en),
.valid_6(PT_L3L4_Plus_TPROJ_FromPlus_L5D4_L3L4_wr_en),
.valid_7(PT_L3L4_Plus_TPROJ_FromPlus_L6D3_L3L4_wr_en),
.valid_8(PT_L3L4_Plus_TPROJ_FromPlus_L6D4_L3L4_wr_en),
.valid_proj_data_stream(PT_L3L4_Plus_To_DataStream_en),
.proj_data_stream(PT_L3L4_Plus_To_DataStream),
.start(start5_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionTransceiver  PT_L5L6_Plus(
.number_in1(TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus_number),
.read_add1(TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus_read_add),
.projin_1(TPROJ_ToPlus_L5D3L6D3_L1_PT_L5L6_Plus),
.number_in2(TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus_number),
.read_add2(TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus_read_add),
.projin_2(TPROJ_ToPlus_L5D3L6D3_L2_PT_L5L6_Plus),
.number_in3(TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus_number),
.read_add3(TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus_read_add),
.projin_3(TPROJ_ToPlus_L5D3L6D3_L3_PT_L5L6_Plus),
.number_in4(TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus_number),
.read_add4(TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus_read_add),
.projin_4(TPROJ_ToPlus_L5D3L6D3_L4_PT_L5L6_Plus),
.number_in5(TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus_number),
.read_add5(TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus_read_add),
.projin_5(TPROJ_ToPlus_L5D3L6D4_L1_PT_L5L6_Plus),
.number_in6(TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus_number),
.read_add6(TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus_read_add),
.projin_6(TPROJ_ToPlus_L5D3L6D4_L2_PT_L5L6_Plus),
.number_in7(TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus_number),
.read_add7(TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus_read_add),
.projin_7(TPROJ_ToPlus_L5D3L6D4_L3_PT_L5L6_Plus),
.number_in8(TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus_number),
.read_add8(TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus_read_add),
.projin_8(TPROJ_ToPlus_L5D3L6D4_L4_PT_L5L6_Plus),
.number_in9(TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus_number),
.read_add9(TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus_read_add),
.projin_9(TPROJ_ToPlus_L5D4L6D4_L1_PT_L5L6_Plus),
.number_in10(TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus_number),
.read_add10(TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus_read_add),
.projin_10(TPROJ_ToPlus_L5D4L6D4_L2_PT_L5L6_Plus),
.number_in11(TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus_number),
.read_add11(TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus_read_add),
.projin_11(TPROJ_ToPlus_L5D4L6D4_L3_PT_L5L6_Plus),
.number_in12(TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus_number),
.read_add12(TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus_read_add),
.projin_12(TPROJ_ToPlus_L5D4L6D4_L4_PT_L5L6_Plus),
.valid_incomming_proj_data_stream(PT_L5L6_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L5L6_Plus_From_DataStream),
.projout_1(PT_L5L6_Plus_TPROJ_FromPlus_L1D3_L5L6),
.projout_2(PT_L5L6_Plus_TPROJ_FromPlus_L1D4_L5L6),
.projout_3(PT_L5L6_Plus_TPROJ_FromPlus_L2D3_L5L6),
.projout_4(PT_L5L6_Plus_TPROJ_FromPlus_L2D4_L5L6),
.projout_5(PT_L5L6_Plus_TPROJ_FromPlus_L3D3_L5L6),
.projout_6(PT_L5L6_Plus_TPROJ_FromPlus_L3D4_L5L6),
.projout_7(PT_L5L6_Plus_TPROJ_FromPlus_L4D3_L5L6),
.projout_8(PT_L5L6_Plus_TPROJ_FromPlus_L4D4_L5L6),
.valid_1(PT_L5L6_Plus_TPROJ_FromPlus_L1D3_L5L6_wr_en),
.valid_2(PT_L5L6_Plus_TPROJ_FromPlus_L1D4_L5L6_wr_en),
.valid_3(PT_L5L6_Plus_TPROJ_FromPlus_L2D3_L5L6_wr_en),
.valid_4(PT_L5L6_Plus_TPROJ_FromPlus_L2D4_L5L6_wr_en),
.valid_5(PT_L5L6_Plus_TPROJ_FromPlus_L3D3_L5L6_wr_en),
.valid_6(PT_L5L6_Plus_TPROJ_FromPlus_L3D4_L5L6_wr_en),
.valid_7(PT_L5L6_Plus_TPROJ_FromPlus_L4D3_L5L6_wr_en),
.valid_8(PT_L5L6_Plus_TPROJ_FromPlus_L4D4_L5L6_wr_en),
.valid_proj_data_stream(PT_L5L6_Plus_To_DataStream_en),
.proj_data_stream(PT_L5L6_Plus_To_DataStream),
.start(start5_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionTransceiver  PT_L1L2_Minus(
.number_in1(TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus_number),
.read_add1(TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus_read_add),
.projin_1(TPROJ_ToMinus_L1D3L2D3_L3_PT_L1L2_Minus),
.number_in2(TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus_number),
.read_add2(TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus_read_add),
.projin_2(TPROJ_ToMinus_L1D3L2D3_L4_PT_L1L2_Minus),
.number_in3(TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus_number),
.read_add3(TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus_read_add),
.projin_3(TPROJ_ToMinus_L1D3L2D3_L5_PT_L1L2_Minus),
.number_in4(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus_number),
.read_add4(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus_read_add),
.projin_4(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L2_Minus),
.number_in5(TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus_number),
.read_add5(TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus_read_add),
.projin_5(TPROJ_ToMinus_L1D3L2D4_L3_PT_L1L2_Minus),
.number_in6(TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus_number),
.read_add6(TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus_read_add),
.projin_6(TPROJ_ToMinus_L1D3L2D4_L4_PT_L1L2_Minus),
.number_in7(TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus_number),
.read_add7(TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus_read_add),
.projin_7(TPROJ_ToMinus_L1D3L2D4_L5_PT_L1L2_Minus),
.number_in8(TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus_number),
.read_add8(TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus_read_add),
.projin_8(TPROJ_ToMinus_L1D3L2D4_L6_PT_L1L2_Minus),
.number_in9(TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus_number),
.read_add9(TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus_read_add),
.projin_9(TPROJ_ToMinus_L1D4L2D4_L3_PT_L1L2_Minus),
.number_in10(TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus_number),
.read_add10(TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus_read_add),
.projin_10(TPROJ_ToMinus_L1D4L2D4_L4_PT_L1L2_Minus),
.number_in11(TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus_number),
.read_add11(TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus_read_add),
.projin_11(TPROJ_ToMinus_L1D4L2D4_L5_PT_L1L2_Minus),
.number_in12(TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus_number),
.read_add12(TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus_read_add),
.projin_12(TPROJ_ToMinus_L1D4L2D4_L6_PT_L1L2_Minus),
.valid_incomming_proj_data_stream(PT_L1L2_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L1L2_Minus_From_DataStream),
.projout_1(PT_L1L2_Minus_TPROJ_FromMinus_L3D3_L1L2),
.projout_2(PT_L1L2_Minus_TPROJ_FromMinus_L3D4_L1L2),
.projout_3(PT_L1L2_Minus_TPROJ_FromMinus_L4D3_L1L2),
.projout_4(PT_L1L2_Minus_TPROJ_FromMinus_L4D4_L1L2),
.projout_5(PT_L1L2_Minus_TPROJ_FromMinus_L5D3_L1L2),
.projout_6(PT_L1L2_Minus_TPROJ_FromMinus_L5D4_L1L2),
.projout_7(PT_L1L2_Minus_TPROJ_FromMinus_L6D3_L1L2),
.projout_8(PT_L1L2_Minus_TPROJ_FromMinus_L6D4_L1L2),
.valid_1(PT_L1L2_Minus_TPROJ_FromMinus_L3D3_L1L2_wr_en),
.valid_2(PT_L1L2_Minus_TPROJ_FromMinus_L3D4_L1L2_wr_en),
.valid_3(PT_L1L2_Minus_TPROJ_FromMinus_L4D3_L1L2_wr_en),
.valid_4(PT_L1L2_Minus_TPROJ_FromMinus_L4D4_L1L2_wr_en),
.valid_5(PT_L1L2_Minus_TPROJ_FromMinus_L5D3_L1L2_wr_en),
.valid_6(PT_L1L2_Minus_TPROJ_FromMinus_L5D4_L1L2_wr_en),
.valid_7(PT_L1L2_Minus_TPROJ_FromMinus_L6D3_L1L2_wr_en),
.valid_8(PT_L1L2_Minus_TPROJ_FromMinus_L6D4_L1L2_wr_en),
.valid_proj_data_stream(PT_L1L2_Minus_To_DataStream_en),
.proj_data_stream(PT_L1L2_Minus_To_DataStream),
.start(start5_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionTransceiver  PT_L3L4_Minus(
.number_in1(TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus_number),
.read_add1(TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus_read_add),
.projin_1(TPROJ_ToMinus_L3D3L4D3_L1_PT_L3L4_Minus),
.number_in2(TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus_number),
.read_add2(TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus_read_add),
.projin_2(TPROJ_ToMinus_L3D3L4D3_L2_PT_L3L4_Minus),
.number_in3(TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus_number),
.read_add3(TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus_read_add),
.projin_3(TPROJ_ToMinus_L3D3L4D3_L5_PT_L3L4_Minus),
.number_in4(TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus_number),
.read_add4(TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus_read_add),
.projin_4(TPROJ_ToMinus_L3D3L4D3_L6_PT_L3L4_Minus),
.number_in5(TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus_number),
.read_add5(TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus_read_add),
.projin_5(TPROJ_ToMinus_L3D3L4D4_L1_PT_L3L4_Minus),
.number_in6(TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus_number),
.read_add6(TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus_read_add),
.projin_6(TPROJ_ToMinus_L3D3L4D4_L2_PT_L3L4_Minus),
.number_in7(TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus_number),
.read_add7(TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus_read_add),
.projin_7(TPROJ_ToMinus_L3D3L4D4_L5_PT_L3L4_Minus),
.number_in8(TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus_number),
.read_add8(TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus_read_add),
.projin_8(TPROJ_ToMinus_L3D3L4D4_L6_PT_L3L4_Minus),
.number_in9(TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus_number),
.read_add9(TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus_read_add),
.projin_9(TPROJ_ToMinus_L3D4L4D4_L1_PT_L3L4_Minus),
.number_in10(TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus_number),
.read_add10(TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus_read_add),
.projin_10(TPROJ_ToMinus_L3D4L4D4_L2_PT_L3L4_Minus),
.number_in11(TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus_number),
.read_add11(TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus_read_add),
.projin_11(TPROJ_ToMinus_L3D4L4D4_L5_PT_L3L4_Minus),
.number_in12(TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus_number),
.read_add12(TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus_read_add),
.projin_12(TPROJ_ToMinus_L3D4L4D4_L6_PT_L3L4_Minus),
.valid_incomming_proj_data_stream(PT_L3L4_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L3L4_Minus_From_DataStream),
.projout_1(PT_L3L4_Minus_TPROJ_FromMinus_L1D3_L3L4),
.projout_2(PT_L3L4_Minus_TPROJ_FromMinus_L1D4_L3L4),
.projout_3(PT_L3L4_Minus_TPROJ_FromMinus_L2D3_L3L4),
.projout_4(PT_L3L4_Minus_TPROJ_FromMinus_L2D4_L3L4),
.projout_5(PT_L3L4_Minus_TPROJ_FromMinus_L5D3_L3L4),
.projout_6(PT_L3L4_Minus_TPROJ_FromMinus_L5D4_L3L4),
.projout_7(PT_L3L4_Minus_TPROJ_FromMinus_L6D3_L3L4),
.projout_8(PT_L3L4_Minus_TPROJ_FromMinus_L6D4_L3L4),
.valid_1(PT_L3L4_Minus_TPROJ_FromMinus_L1D3_L3L4_wr_en),
.valid_2(PT_L3L4_Minus_TPROJ_FromMinus_L1D4_L3L4_wr_en),
.valid_3(PT_L3L4_Minus_TPROJ_FromMinus_L2D3_L3L4_wr_en),
.valid_4(PT_L3L4_Minus_TPROJ_FromMinus_L2D4_L3L4_wr_en),
.valid_5(PT_L3L4_Minus_TPROJ_FromMinus_L5D3_L3L4_wr_en),
.valid_6(PT_L3L4_Minus_TPROJ_FromMinus_L5D4_L3L4_wr_en),
.valid_7(PT_L3L4_Minus_TPROJ_FromMinus_L6D3_L3L4_wr_en),
.valid_8(PT_L3L4_Minus_TPROJ_FromMinus_L6D4_L3L4_wr_en),
.valid_proj_data_stream(PT_L3L4_Minus_To_DataStream_en),
.proj_data_stream(PT_L3L4_Minus_To_DataStream),
.start(start5_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionTransceiver  PT_L5L6_Minus(
.number_in1(TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus_number),
.read_add1(TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus_read_add),
.projin_1(TPROJ_ToMinus_L5D3L6D3_L1_PT_L5L6_Minus),
.number_in2(TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus_number),
.read_add2(TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus_read_add),
.projin_2(TPROJ_ToMinus_L5D3L6D3_L2_PT_L5L6_Minus),
.number_in3(TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus_number),
.read_add3(TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus_read_add),
.projin_3(TPROJ_ToMinus_L5D3L6D3_L3_PT_L5L6_Minus),
.number_in4(TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus_number),
.read_add4(TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus_read_add),
.projin_4(TPROJ_ToMinus_L5D3L6D3_L4_PT_L5L6_Minus),
.number_in5(TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus_number),
.read_add5(TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus_read_add),
.projin_5(TPROJ_ToMinus_L5D3L6D4_L1_PT_L5L6_Minus),
.number_in6(TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus_number),
.read_add6(TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus_read_add),
.projin_6(TPROJ_ToMinus_L5D3L6D4_L2_PT_L5L6_Minus),
.number_in7(TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus_number),
.read_add7(TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus_read_add),
.projin_7(TPROJ_ToMinus_L5D3L6D4_L3_PT_L5L6_Minus),
.number_in8(TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus_number),
.read_add8(TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus_read_add),
.projin_8(TPROJ_ToMinus_L5D3L6D4_L4_PT_L5L6_Minus),
.number_in9(TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus_number),
.read_add9(TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus_read_add),
.projin_9(TPROJ_ToMinus_L5D4L6D4_L1_PT_L5L6_Minus),
.number_in10(TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus_number),
.read_add10(TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus_read_add),
.projin_10(TPROJ_ToMinus_L5D4L6D4_L2_PT_L5L6_Minus),
.number_in11(TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus_number),
.read_add11(TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus_read_add),
.projin_11(TPROJ_ToMinus_L5D4L6D4_L3_PT_L5L6_Minus),
.number_in12(TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus_number),
.read_add12(TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus_read_add),
.projin_12(TPROJ_ToMinus_L5D4L6D4_L4_PT_L5L6_Minus),
.valid_incomming_proj_data_stream(PT_L5L6_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L5L6_Minus_From_DataStream),
.projout_1(PT_L5L6_Minus_TPROJ_FromMinus_L1D3_L5L6),
.projout_2(PT_L5L6_Minus_TPROJ_FromMinus_L1D4_L5L6),
.projout_3(PT_L5L6_Minus_TPROJ_FromMinus_L2D3_L5L6),
.projout_4(PT_L5L6_Minus_TPROJ_FromMinus_L2D4_L5L6),
.projout_5(PT_L5L6_Minus_TPROJ_FromMinus_L3D3_L5L6),
.projout_6(PT_L5L6_Minus_TPROJ_FromMinus_L3D4_L5L6),
.projout_7(PT_L5L6_Minus_TPROJ_FromMinus_L4D3_L5L6),
.projout_8(PT_L5L6_Minus_TPROJ_FromMinus_L4D4_L5L6),
.valid_1(PT_L5L6_Minus_TPROJ_FromMinus_L1D3_L5L6_wr_en),
.valid_2(PT_L5L6_Minus_TPROJ_FromMinus_L1D4_L5L6_wr_en),
.valid_3(PT_L5L6_Minus_TPROJ_FromMinus_L2D3_L5L6_wr_en),
.valid_4(PT_L5L6_Minus_TPROJ_FromMinus_L2D4_L5L6_wr_en),
.valid_5(PT_L5L6_Minus_TPROJ_FromMinus_L3D3_L5L6_wr_en),
.valid_6(PT_L5L6_Minus_TPROJ_FromMinus_L3D4_L5L6_wr_en),
.valid_7(PT_L5L6_Minus_TPROJ_FromMinus_L4D3_L5L6_wr_en),
.valid_8(PT_L5L6_Minus_TPROJ_FromMinus_L4D4_L5L6_wr_en),
.valid_proj_data_stream(PT_L5L6_Minus_To_DataStream_en),
.proj_data_stream(PT_L5L6_Minus_To_DataStream),
.start(start5_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b1) PR_L1D3_L3L4(
.number_in1(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_number),
.read_add1(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4),
.number_in2(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_number),
.read_add2(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4),
.number_in3(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_number),
.read_add3(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4),
.number_in4(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_number),
.read_add4(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4),
.number_in5(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_number),
.read_add5(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4),
.vmprojoutPHI1Z1(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z2),
.allprojout(PR_L1D3_L3L4_AP_L3L4_L1D3),
.valid_data(PR_L1D3_L3L4_AP_L3L4_L1D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3Z2_wr_en),
.start(start6_5),
.done(done6_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b1) PR_L1D4_L3L4(
.number_in1(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_number),
.read_add1(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4),
.number_in2(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_number),
.read_add2(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4),
.number_in3(TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4_number),
.read_add3(TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L1D4_PR_L1D4_L3L4),
.number_in4(TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4_number),
.read_add4(TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L1D4_PR_L1D4_L3L4),
.number_in5(TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4_number),
.read_add5(TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L1D4_PR_L1D4_L3L4),
.vmprojoutPHI1Z1(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z2),
.allprojout(PR_L1D4_L3L4_AP_L3L4_L1D4),
.valid_data(PR_L1D4_L3L4_AP_L3L4_L1D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b1) PR_L2D3_L3L4(
.number_in1(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_number),
.read_add1(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4),
.number_in2(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_number),
.read_add2(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4),
.number_in3(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_number),
.read_add3(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4),
.number_in4(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_number),
.read_add4(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4),
.number_in5(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_number),
.read_add5(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4),
.vmprojoutPHI1Z1(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z2),
.vmprojoutPHI4Z1(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z1),
.vmprojoutPHI4Z2(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z2),
.allprojout(PR_L2D3_L3L4_AP_L3L4_L2D3),
.valid_data(PR_L2D3_L3L4_AP_L3L4_L2D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b1) PR_L2D4_L3L4(
.number_in1(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_number),
.read_add1(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4),
.number_in2(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_number),
.read_add2(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4),
.number_in3(TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4_number),
.read_add3(TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L2D4_PR_L2D4_L3L4),
.number_in4(TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4_number),
.read_add4(TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L2D4_PR_L2D4_L3L4),
.number_in5(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_number),
.read_add5(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4),
.vmprojoutPHI1Z1(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z2),
.vmprojoutPHI4Z1(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z1),
.vmprojoutPHI4Z2(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z2),
.allprojout(PR_L2D4_L3L4_AP_L3L4_L2D4),
.valid_data(PR_L2D4_L3L4_AP_L3L4_L2D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b0) PR_L5D3_L3L4(
.number_in1(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_number),
.read_add1(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4),
.number_in2(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_number),
.read_add2(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4),
.number_in3(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_number),
.read_add3(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4),
.number_in4(TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4_number),
.read_add4(TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L5D3_PR_L5D3_L3L4),
.number_in5(TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4_number),
.read_add5(TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L5D3_PR_L5D3_L3L4),
.vmprojoutPHI1Z1(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z2),
.allprojout(PR_L5D3_L3L4_AP_L3L4_L5D3),
.valid_data(PR_L5D3_L3L4_AP_L3L4_L5D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b0) PR_L5D4_L3L4(
.number_in1(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_number),
.read_add1(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4),
.number_in2(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_number),
.read_add2(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4),
.number_in3(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_number),
.read_add3(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4),
.number_in4(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_number),
.read_add4(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4),
.number_in5(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_number),
.read_add5(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4),
.vmprojoutPHI1Z1(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z2),
.allprojout(PR_L5D4_L3L4_AP_L3L4_L5D4),
.valid_data(PR_L5D4_L3L4_AP_L3L4_L5D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b0) PR_L6D3_L3L4(
.number_in1(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_number),
.read_add1(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4),
.number_in2(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_number),
.read_add2(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4),
.number_in3(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_number),
.read_add3(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4),
.number_in4(TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4_number),
.read_add4(TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L6D3_PR_L6D3_L3L4),
.number_in5(TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4_number),
.read_add5(TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L6D3_PR_L6D3_L3L4),
.vmprojoutPHI1Z1(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z2),
.vmprojoutPHI4Z1(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z1),
.vmprojoutPHI4Z2(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z2),
.allprojout(PR_L6D3_L3L4_AP_L3L4_L6D3),
.valid_data(PR_L6D3_L3L4_AP_L3L4_L6D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b0) PR_L6D4_L3L4(
.number_in1(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_number),
.read_add1(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4),
.number_in2(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_number),
.read_add2(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4),
.number_in3(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_number),
.read_add3(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4),
.number_in4(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_number),
.read_add4(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4),
.number_in5(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_number),
.read_add5(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4),
.vmprojoutPHI1Z1(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z2),
.vmprojoutPHI4Z1(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z1),
.vmprojoutPHI4Z2(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z2),
.allprojout(PR_L6D4_L3L4_AP_L3L4_L6D4),
.valid_data(PR_L6D4_L3L4_AP_L3L4_L6D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b1) PR_L3D3_L1L2(
.number_in1(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_number),
.read_add1(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2),
.number_in2(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_number),
.read_add2(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2),
.number_in3(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_number),
.read_add3(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2),
.number_in4(TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2_number),
.read_add4(TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L3D3_PR_L3D3_L1L2),
.number_in5(TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2_number),
.read_add5(TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L3D3_PR_L3D3_L1L2),
.vmprojoutPHI1Z1(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z2),
.allprojout(PR_L3D3_L1L2_AP_L1L2_L3D3),
.valid_data(PR_L3D3_L1L2_AP_L1L2_L3D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b1) PR_L3D4_L1L2(
.number_in1(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_number),
.read_add1(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2),
.number_in2(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_number),
.read_add2(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2),
.number_in3(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_number),
.read_add3(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2),
.number_in4(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_number),
.read_add4(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2),
.number_in5(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_number),
.read_add5(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2),
.vmprojoutPHI1Z1(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z2),
.allprojout(PR_L3D4_L1L2_AP_L1L2_L3D4),
.valid_data(PR_L3D4_L1L2_AP_L1L2_L3D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b0) PR_L4D3_L1L2(
.number_in1(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_number),
.read_add1(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2),
.number_in2(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_number),
.read_add2(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2),
.number_in3(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_number),
.read_add3(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2),
.number_in4(TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2_number),
.read_add4(TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L4D3_PR_L4D3_L1L2),
.number_in5(TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2_number),
.read_add5(TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L4D3_PR_L4D3_L1L2),
.vmprojoutPHI1Z1(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z2),
.vmprojoutPHI4Z1(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z1),
.vmprojoutPHI4Z2(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z2),
.allprojout(PR_L4D3_L1L2_AP_L1L2_L4D3),
.valid_data(PR_L4D3_L1L2_AP_L1L2_L4D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b0) PR_L4D4_L1L2(
.number_in1(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_number),
.read_add1(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2),
.number_in2(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_number),
.read_add2(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2),
.number_in3(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_number),
.read_add3(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2),
.number_in4(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_number),
.read_add4(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2),
.number_in5(TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2_number),
.read_add5(TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L4D4_PR_L4D4_L1L2),
.vmprojoutPHI1Z1(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z2),
.vmprojoutPHI4Z1(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z1),
.vmprojoutPHI4Z2(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z2),
.allprojout(PR_L4D4_L1L2_AP_L1L2_L4D4),
.valid_data(PR_L4D4_L1L2_AP_L1L2_L4D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b0) PR_L5D3_L1L2(
.number_in1(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_number),
.read_add1(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2),
.number_in2(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_number),
.read_add2(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2),
.number_in3(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_number),
.read_add3(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2),
.number_in4(TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2_number),
.read_add4(TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L5D3_PR_L5D3_L1L2),
.number_in5(TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2_number),
.read_add5(TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L5D3_PR_L5D3_L1L2),
.vmprojoutPHI1Z1(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z2),
.allprojout(PR_L5D3_L1L2_AP_L1L2_L5D3),
.valid_data(PR_L5D3_L1L2_AP_L1L2_L5D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b0) PR_L5D4_L1L2(
.number_in1(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_number),
.read_add1(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2),
.number_in2(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_number),
.read_add2(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2),
.number_in3(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_number),
.read_add3(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2),
.number_in4(TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2_number),
.read_add4(TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L5D4_PR_L5D4_L1L2),
.number_in5(TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2_number),
.read_add5(TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L5D4_PR_L5D4_L1L2),
.vmprojoutPHI1Z1(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z2),
.allprojout(PR_L5D4_L1L2_AP_L1L2_L5D4),
.valid_data(PR_L5D4_L1L2_AP_L1L2_L5D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b0) PR_L6D3_L1L2(
.number_in1(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_number),
.read_add1(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2),
.number_in2(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_number),
.read_add2(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2),
.number_in3(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_number),
.read_add3(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2),
.number_in4(TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2_number),
.read_add4(TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L6D3_PR_L6D3_L1L2),
.number_in5(TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2_number),
.read_add5(TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L6D3_PR_L6D3_L1L2),
.vmprojoutPHI1Z1(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z2),
.vmprojoutPHI4Z1(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z1),
.vmprojoutPHI4Z2(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z2),
.allprojout(PR_L6D3_L1L2_AP_L1L2_L6D3),
.valid_data(PR_L6D3_L1L2_AP_L1L2_L6D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b0) PR_L6D4_L1L2(
.number_in1(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_number),
.read_add1(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2),
.number_in2(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_number),
.read_add2(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2),
.number_in3(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_number),
.read_add3(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2),
.number_in4(TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2_number),
.read_add4(TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L6D4_PR_L6D4_L1L2),
.number_in5(TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2_number),
.read_add5(TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L6D4_PR_L6D4_L1L2),
.vmprojoutPHI1Z1(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z2),
.vmprojoutPHI4Z1(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z1),
.vmprojoutPHI4Z2(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z2),
.allprojout(PR_L6D4_L1L2_AP_L1L2_L6D4),
.valid_data(PR_L6D4_L1L2_AP_L1L2_L6D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b1) PR_L1D3_L5L6(
.number_in1(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_number),
.read_add1(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6),
.number_in2(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_number),
.read_add2(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6),
.number_in3(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_number),
.read_add3(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6),
.number_in4(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_number),
.read_add4(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6),
.number_in5(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_number),
.read_add5(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6),
.vmprojoutPHI1Z1(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z2),
.allprojout(PR_L1D3_L5L6_AP_L5L6_L1D3),
.valid_data(PR_L1D3_L5L6_AP_L5L6_L1D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b1) PR_L1D4_L5L6(
.number_in1(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_number),
.read_add1(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6),
.number_in2(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_number),
.read_add2(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6),
.number_in3(TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6_number),
.read_add3(TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L1D4_PR_L1D4_L5L6),
.number_in4(TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6_number),
.read_add4(TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L1D4_PR_L1D4_L5L6),
.number_in5(TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6_number),
.read_add5(TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L1D4_PR_L1D4_L5L6),
.vmprojoutPHI1Z1(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z2),
.allprojout(PR_L1D4_L5L6_AP_L5L6_L1D4),
.valid_data(PR_L1D4_L5L6_AP_L5L6_L1D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b1) PR_L2D3_L5L6(
.number_in1(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_number),
.read_add1(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6),
.number_in2(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_number),
.read_add2(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6),
.number_in3(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_number),
.read_add3(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6),
.number_in4(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_number),
.read_add4(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6),
.number_in5(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_number),
.read_add5(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6),
.vmprojoutPHI1Z1(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z2),
.vmprojoutPHI4Z1(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z1),
.vmprojoutPHI4Z2(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z2),
.allprojout(PR_L2D3_L5L6_AP_L5L6_L2D3),
.valid_data(PR_L2D3_L5L6_AP_L5L6_L2D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b1) PR_L2D4_L5L6(
.number_in1(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_number),
.read_add1(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6),
.number_in2(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_number),
.read_add2(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6),
.number_in3(TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6_number),
.read_add3(TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L2D4_PR_L2D4_L5L6),
.number_in4(TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6_number),
.read_add4(TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L2D4_PR_L2D4_L5L6),
.number_in5(TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6_number),
.read_add5(TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L2D4_PR_L2D4_L5L6),
.vmprojoutPHI1Z1(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z2),
.vmprojoutPHI4Z1(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z1),
.vmprojoutPHI4Z2(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z2),
.allprojout(PR_L2D4_L5L6_AP_L5L6_L2D4),
.valid_data(PR_L2D4_L5L6_AP_L5L6_L2D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b1) PR_L3D3_L5L6(
.number_in1(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_number),
.read_add1(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6),
.number_in2(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_number),
.read_add2(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6),
.number_in3(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_number),
.read_add3(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6),
.number_in4(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_number),
.read_add4(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6),
.number_in5(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_number),
.read_add5(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6),
.vmprojoutPHI1Z1(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z2),
.allprojout(PR_L3D3_L5L6_AP_L5L6_L3D3),
.valid_data(PR_L3D3_L5L6_AP_L5L6_L3D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b1,1'b1) PR_L3D4_L5L6(
.number_in1(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_number),
.read_add1(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6),
.number_in2(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_number),
.read_add2(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6),
.number_in3(TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6_number),
.read_add3(TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L3D4_PR_L3D4_L5L6),
.number_in4(TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6_number),
.read_add4(TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L3D4_PR_L3D4_L5L6),
.number_in5(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_number),
.read_add5(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6),
.vmprojoutPHI1Z1(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z2),
.allprojout(PR_L3D4_L5L6_AP_L5L6_L3D4),
.valid_data(PR_L3D4_L5L6_AP_L5L6_L3D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b0) PR_L4D3_L5L6(
.number_in1(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_number),
.read_add1(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6),
.number_in2(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_number),
.read_add2(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6),
.number_in3(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_number),
.read_add3(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6),
.number_in4(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_number),
.read_add4(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6),
.number_in5(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_number),
.read_add5(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6),
.vmprojoutPHI1Z1(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z1),
.vmprojoutPHI1Z2(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z2),
.vmprojoutPHI2Z1(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z1),
.vmprojoutPHI2Z2(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z2),
.vmprojoutPHI3Z1(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z1),
.vmprojoutPHI3Z2(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z2),
.vmprojoutPHI4Z1(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z1),
.vmprojoutPHI4Z2(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z2),
.allprojout(PR_L4D3_L5L6_AP_L5L6_L4D3),
.valid_data(PR_L4D3_L5L6_AP_L5L6_L4D3_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


ProjectionRouter #(1'b0,1'b0) PR_L4D4_L5L6(
.number_in1(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_number),
.read_add1(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6),
.number_in2(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_number),
.read_add2(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6),
.number_in3(TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6_number),
.read_add3(TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L4D4_PR_L4D4_L5L6),
.number_in4(TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6_number),
.read_add4(TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L4D4_PR_L4D4_L5L6),
.number_in5(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_number),
.read_add5(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6),
.vmprojoutPHI1Z1(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z1),
.vmprojoutPHI1Z2(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z2),
.vmprojoutPHI2Z1(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z1),
.vmprojoutPHI2Z2(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z2),
.vmprojoutPHI3Z1(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z1),
.vmprojoutPHI3Z2(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z2),
.vmprojoutPHI4Z1(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z1),
.vmprojoutPHI4Z2(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z2),
.allprojout(PR_L4D4_L5L6_AP_L5L6_L4D4),
.valid_data(PR_L4D4_L5L6_AP_L5L6_L4D4_wr_en),
.vmprojoutPHI1Z1_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z1_wr_en),
.vmprojoutPHI1Z2_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1Z2_wr_en),
.vmprojoutPHI2Z1_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z1_wr_en),
.vmprojoutPHI2Z2_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2Z2_wr_en),
.vmprojoutPHI3Z1_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z1_wr_en),
.vmprojoutPHI3Z2_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3Z2_wr_en),
.vmprojoutPHI4Z1_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z1_wr_en),
.vmprojoutPHI4Z2_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4Z2_wr_en),
.start(start6_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D3PHI1Z1(
.number_in1(VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1_number),
.read_add1(VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1_read_add),
.vmstubin(VMS_L1D3PHI1Z1n7_ME_L3L4_L1D3PHI1Z1),
.number_in2(VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1_number),
.read_add2(VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI1Z1_ME_L3L4_L1D3PHI1Z1),
.matchout(ME_L3L4_L1D3PHI1Z1_CM_L3L4_L1D3PHI1Z1),
.valid_data(ME_L3L4_L1D3PHI1Z1_CM_L3L4_L1D3PHI1Z1_wr_en),
.start(start7_5),
.done(done7_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D3PHI1Z2(
.number_in1(VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2_number),
.read_add1(VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2_read_add),
.vmstubin(VMS_L1D3PHI1Z2n7_ME_L3L4_L1D3PHI1Z2),
.number_in2(VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2_number),
.read_add2(VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI1Z2_ME_L3L4_L1D3PHI1Z2),
.matchout(ME_L3L4_L1D3PHI1Z2_CM_L3L4_L1D3PHI1Z2),
.valid_data(ME_L3L4_L1D3PHI1Z2_CM_L3L4_L1D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D3PHI2Z1(
.number_in1(VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1_number),
.read_add1(VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1_read_add),
.vmstubin(VMS_L1D3PHI2Z1n7_ME_L3L4_L1D3PHI2Z1),
.number_in2(VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1_number),
.read_add2(VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI2Z1_ME_L3L4_L1D3PHI2Z1),
.matchout(ME_L3L4_L1D3PHI2Z1_CM_L3L4_L1D3PHI2Z1),
.valid_data(ME_L3L4_L1D3PHI2Z1_CM_L3L4_L1D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D3PHI2Z2(
.number_in1(VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2_number),
.read_add1(VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2_read_add),
.vmstubin(VMS_L1D3PHI2Z2n7_ME_L3L4_L1D3PHI2Z2),
.number_in2(VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2_number),
.read_add2(VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI2Z2_ME_L3L4_L1D3PHI2Z2),
.matchout(ME_L3L4_L1D3PHI2Z2_CM_L3L4_L1D3PHI2Z2),
.valid_data(ME_L3L4_L1D3PHI2Z2_CM_L3L4_L1D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D3PHI3Z1(
.number_in1(VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1_number),
.read_add1(VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1_read_add),
.vmstubin(VMS_L1D3PHI3Z1n7_ME_L3L4_L1D3PHI3Z1),
.number_in2(VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1_number),
.read_add2(VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI3Z1_ME_L3L4_L1D3PHI3Z1),
.matchout(ME_L3L4_L1D3PHI3Z1_CM_L3L4_L1D3PHI3Z1),
.valid_data(ME_L3L4_L1D3PHI3Z1_CM_L3L4_L1D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D3PHI3Z2(
.number_in1(VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2_number),
.read_add1(VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2_read_add),
.vmstubin(VMS_L1D3PHI3Z2n7_ME_L3L4_L1D3PHI3Z2),
.number_in2(VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2_number),
.read_add2(VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI3Z2_ME_L3L4_L1D3PHI3Z2),
.matchout(ME_L3L4_L1D3PHI3Z2_CM_L3L4_L1D3PHI3Z2),
.valid_data(ME_L3L4_L1D3PHI3Z2_CM_L3L4_L1D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D4PHI1Z1(
.number_in1(VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1_number),
.read_add1(VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1_read_add),
.vmstubin(VMS_L1D4PHI1Z1n3_ME_L3L4_L1D4PHI1Z1),
.number_in2(VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1_number),
.read_add2(VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI1Z1_ME_L3L4_L1D4PHI1Z1),
.matchout(ME_L3L4_L1D4PHI1Z1_CM_L3L4_L1D4PHI1Z1),
.valid_data(ME_L3L4_L1D4PHI1Z1_CM_L3L4_L1D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D4PHI1Z2(
.number_in1(VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2_number),
.read_add1(VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI1Z2_ME_L3L4_L1D4PHI1Z2),
.number_in2(VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2_number),
.read_add2(VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2_read_add),
.vmstubin(VMS_L1D4PHI1Z2n1_ME_L3L4_L1D4PHI1Z2),
.matchout(ME_L3L4_L1D4PHI1Z2_CM_L3L4_L1D4PHI1Z2),
.valid_data(ME_L3L4_L1D4PHI1Z2_CM_L3L4_L1D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D4PHI2Z1(
.number_in1(VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1_number),
.read_add1(VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1_read_add),
.vmstubin(VMS_L1D4PHI2Z1n3_ME_L3L4_L1D4PHI2Z1),
.number_in2(VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1_number),
.read_add2(VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI2Z1_ME_L3L4_L1D4PHI2Z1),
.matchout(ME_L3L4_L1D4PHI2Z1_CM_L3L4_L1D4PHI2Z1),
.valid_data(ME_L3L4_L1D4PHI2Z1_CM_L3L4_L1D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D4PHI2Z2(
.number_in1(VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2_number),
.read_add1(VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI2Z2_ME_L3L4_L1D4PHI2Z2),
.number_in2(VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2_number),
.read_add2(VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2_read_add),
.vmstubin(VMS_L1D4PHI2Z2n1_ME_L3L4_L1D4PHI2Z2),
.matchout(ME_L3L4_L1D4PHI2Z2_CM_L3L4_L1D4PHI2Z2),
.valid_data(ME_L3L4_L1D4PHI2Z2_CM_L3L4_L1D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D4PHI3Z1(
.number_in1(VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1_number),
.read_add1(VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1_read_add),
.vmstubin(VMS_L1D4PHI3Z1n3_ME_L3L4_L1D4PHI3Z1),
.number_in2(VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1_number),
.read_add2(VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI3Z1_ME_L3L4_L1D4PHI3Z1),
.matchout(ME_L3L4_L1D4PHI3Z1_CM_L3L4_L1D4PHI3Z1),
.valid_data(ME_L3L4_L1D4PHI3Z1_CM_L3L4_L1D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L1D4PHI3Z2(
.number_in1(VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2_number),
.read_add1(VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI3Z2_ME_L3L4_L1D4PHI3Z2),
.number_in2(VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2_number),
.read_add2(VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2_read_add),
.vmstubin(VMS_L1D4PHI3Z2n1_ME_L3L4_L1D4PHI3Z2),
.matchout(ME_L3L4_L1D4PHI3Z2_CM_L3L4_L1D4PHI3Z2),
.valid_data(ME_L3L4_L1D4PHI3Z2_CM_L3L4_L1D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D3PHI1Z1(
.number_in1(VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1_number),
.read_add1(VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1_read_add),
.vmstubin(VMS_L2D3PHI1Z1n2_ME_L3L4_L2D3PHI1Z1),
.number_in2(VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1_number),
.read_add2(VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI1Z1_ME_L3L4_L2D3PHI1Z1),
.matchout(ME_L3L4_L2D3PHI1Z1_CM_L3L4_L2D3PHI1Z1),
.valid_data(ME_L3L4_L2D3PHI1Z1_CM_L3L4_L2D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D3PHI1Z2(
.number_in1(VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2_number),
.read_add1(VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2_read_add),
.vmstubin(VMS_L2D3PHI1Z2n3_ME_L3L4_L2D3PHI1Z2),
.number_in2(VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2_number),
.read_add2(VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI1Z2_ME_L3L4_L2D3PHI1Z2),
.matchout(ME_L3L4_L2D3PHI1Z2_CM_L3L4_L2D3PHI1Z2),
.valid_data(ME_L3L4_L2D3PHI1Z2_CM_L3L4_L2D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D3PHI2Z1(
.number_in1(VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1_number),
.read_add1(VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1_read_add),
.vmstubin(VMS_L2D3PHI2Z1n3_ME_L3L4_L2D3PHI2Z1),
.number_in2(VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1_number),
.read_add2(VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI2Z1_ME_L3L4_L2D3PHI2Z1),
.matchout(ME_L3L4_L2D3PHI2Z1_CM_L3L4_L2D3PHI2Z1),
.valid_data(ME_L3L4_L2D3PHI2Z1_CM_L3L4_L2D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D3PHI2Z2(
.number_in1(VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2_number),
.read_add1(VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2_read_add),
.vmstubin(VMS_L2D3PHI2Z2n5_ME_L3L4_L2D3PHI2Z2),
.number_in2(VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2_number),
.read_add2(VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI2Z2_ME_L3L4_L2D3PHI2Z2),
.matchout(ME_L3L4_L2D3PHI2Z2_CM_L3L4_L2D3PHI2Z2),
.valid_data(ME_L3L4_L2D3PHI2Z2_CM_L3L4_L2D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D3PHI3Z1(
.number_in1(VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1_number),
.read_add1(VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1_read_add),
.vmstubin(VMS_L2D3PHI3Z1n3_ME_L3L4_L2D3PHI3Z1),
.number_in2(VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1_number),
.read_add2(VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI3Z1_ME_L3L4_L2D3PHI3Z1),
.matchout(ME_L3L4_L2D3PHI3Z1_CM_L3L4_L2D3PHI3Z1),
.valid_data(ME_L3L4_L2D3PHI3Z1_CM_L3L4_L2D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D3PHI3Z2(
.number_in1(VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2_number),
.read_add1(VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2_read_add),
.vmstubin(VMS_L2D3PHI3Z2n5_ME_L3L4_L2D3PHI3Z2),
.number_in2(VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2_number),
.read_add2(VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI3Z2_ME_L3L4_L2D3PHI3Z2),
.matchout(ME_L3L4_L2D3PHI3Z2_CM_L3L4_L2D3PHI3Z2),
.valid_data(ME_L3L4_L2D3PHI3Z2_CM_L3L4_L2D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D3PHI4Z1(
.number_in1(VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1_number),
.read_add1(VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1_read_add),
.vmstubin(VMS_L2D3PHI4Z1n2_ME_L3L4_L2D3PHI4Z1),
.number_in2(VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1_number),
.read_add2(VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI4Z1_ME_L3L4_L2D3PHI4Z1),
.matchout(ME_L3L4_L2D3PHI4Z1_CM_L3L4_L2D3PHI4Z1),
.valid_data(ME_L3L4_L2D3PHI4Z1_CM_L3L4_L2D3PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D3PHI4Z2(
.number_in1(VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2_number),
.read_add1(VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2_read_add),
.vmstubin(VMS_L2D3PHI4Z2n3_ME_L3L4_L2D3PHI4Z2),
.number_in2(VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2_number),
.read_add2(VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI4Z2_ME_L3L4_L2D3PHI4Z2),
.matchout(ME_L3L4_L2D3PHI4Z2_CM_L3L4_L2D3PHI4Z2),
.valid_data(ME_L3L4_L2D3PHI4Z2_CM_L3L4_L2D3PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D4PHI1Z1(
.number_in1(VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1_number),
.read_add1(VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1_read_add),
.vmstubin(VMS_L2D4PHI1Z1n3_ME_L3L4_L2D4PHI1Z1),
.number_in2(VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1_number),
.read_add2(VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI1Z1_ME_L3L4_L2D4PHI1Z1),
.matchout(ME_L3L4_L2D4PHI1Z1_CM_L3L4_L2D4PHI1Z1),
.valid_data(ME_L3L4_L2D4PHI1Z1_CM_L3L4_L2D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D4PHI1Z2(
.number_in1(VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2_number),
.read_add1(VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2_read_add),
.vmstubin(VMS_L2D4PHI1Z2n3_ME_L3L4_L2D4PHI1Z2),
.number_in2(VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2_number),
.read_add2(VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI1Z2_ME_L3L4_L2D4PHI1Z2),
.matchout(ME_L3L4_L2D4PHI1Z2_CM_L3L4_L2D4PHI1Z2),
.valid_data(ME_L3L4_L2D4PHI1Z2_CM_L3L4_L2D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D4PHI2Z1(
.number_in1(VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1_number),
.read_add1(VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1_read_add),
.vmstubin(VMS_L2D4PHI2Z1n5_ME_L3L4_L2D4PHI2Z1),
.number_in2(VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1_number),
.read_add2(VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI2Z1_ME_L3L4_L2D4PHI2Z1),
.matchout(ME_L3L4_L2D4PHI2Z1_CM_L3L4_L2D4PHI2Z1),
.valid_data(ME_L3L4_L2D4PHI2Z1_CM_L3L4_L2D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D4PHI2Z2(
.number_in1(VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2_number),
.read_add1(VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2_read_add),
.vmstubin(VMS_L2D4PHI2Z2n5_ME_L3L4_L2D4PHI2Z2),
.number_in2(VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2_number),
.read_add2(VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI2Z2_ME_L3L4_L2D4PHI2Z2),
.matchout(ME_L3L4_L2D4PHI2Z2_CM_L3L4_L2D4PHI2Z2),
.valid_data(ME_L3L4_L2D4PHI2Z2_CM_L3L4_L2D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D4PHI3Z1(
.number_in1(VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1_number),
.read_add1(VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1_read_add),
.vmstubin(VMS_L2D4PHI3Z1n5_ME_L3L4_L2D4PHI3Z1),
.number_in2(VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1_number),
.read_add2(VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI3Z1_ME_L3L4_L2D4PHI3Z1),
.matchout(ME_L3L4_L2D4PHI3Z1_CM_L3L4_L2D4PHI3Z1),
.valid_data(ME_L3L4_L2D4PHI3Z1_CM_L3L4_L2D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D4PHI3Z2(
.number_in1(VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2_number),
.read_add1(VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2_read_add),
.vmstubin(VMS_L2D4PHI3Z2n5_ME_L3L4_L2D4PHI3Z2),
.number_in2(VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2_number),
.read_add2(VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI3Z2_ME_L3L4_L2D4PHI3Z2),
.matchout(ME_L3L4_L2D4PHI3Z2_CM_L3L4_L2D4PHI3Z2),
.valid_data(ME_L3L4_L2D4PHI3Z2_CM_L3L4_L2D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D4PHI4Z1(
.number_in1(VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1_number),
.read_add1(VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1_read_add),
.vmstubin(VMS_L2D4PHI4Z1n3_ME_L3L4_L2D4PHI4Z1),
.number_in2(VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1_number),
.read_add2(VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI4Z1_ME_L3L4_L2D4PHI4Z1),
.matchout(ME_L3L4_L2D4PHI4Z1_CM_L3L4_L2D4PHI4Z1),
.valid_data(ME_L3L4_L2D4PHI4Z1_CM_L3L4_L2D4PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L2D4PHI4Z2(
.number_in1(VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2_number),
.read_add1(VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2_read_add),
.vmstubin(VMS_L2D4PHI4Z2n3_ME_L3L4_L2D4PHI4Z2),
.number_in2(VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2_number),
.read_add2(VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI4Z2_ME_L3L4_L2D4PHI4Z2),
.matchout(ME_L3L4_L2D4PHI4Z2_CM_L3L4_L2D4PHI4Z2),
.valid_data(ME_L3L4_L2D4PHI4Z2_CM_L3L4_L2D4PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D3PHI1Z1(
.number_in1(VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1_number),
.read_add1(VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1_read_add),
.vmstubin(VMS_L5D3PHI1Z1n5_ME_L3L4_L5D3PHI1Z1),
.number_in2(VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1_number),
.read_add2(VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI1Z1_ME_L3L4_L5D3PHI1Z1),
.matchout(ME_L3L4_L5D3PHI1Z1_CM_L3L4_L5D3PHI1Z1),
.valid_data(ME_L3L4_L5D3PHI1Z1_CM_L3L4_L5D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D3PHI1Z2(
.number_in1(VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2_number),
.read_add1(VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2_read_add),
.vmstubin(VMS_L5D3PHI1Z2n5_ME_L3L4_L5D3PHI1Z2),
.number_in2(VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2_number),
.read_add2(VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI1Z2_ME_L3L4_L5D3PHI1Z2),
.matchout(ME_L3L4_L5D3PHI1Z2_CM_L3L4_L5D3PHI1Z2),
.valid_data(ME_L3L4_L5D3PHI1Z2_CM_L3L4_L5D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D3PHI2Z1(
.number_in1(VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1_number),
.read_add1(VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1_read_add),
.vmstubin(VMS_L5D3PHI2Z1n5_ME_L3L4_L5D3PHI2Z1),
.number_in2(VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1_number),
.read_add2(VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI2Z1_ME_L3L4_L5D3PHI2Z1),
.matchout(ME_L3L4_L5D3PHI2Z1_CM_L3L4_L5D3PHI2Z1),
.valid_data(ME_L3L4_L5D3PHI2Z1_CM_L3L4_L5D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D3PHI2Z2(
.number_in1(VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2_number),
.read_add1(VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2_read_add),
.vmstubin(VMS_L5D3PHI2Z2n5_ME_L3L4_L5D3PHI2Z2),
.number_in2(VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2_number),
.read_add2(VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI2Z2_ME_L3L4_L5D3PHI2Z2),
.matchout(ME_L3L4_L5D3PHI2Z2_CM_L3L4_L5D3PHI2Z2),
.valid_data(ME_L3L4_L5D3PHI2Z2_CM_L3L4_L5D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D3PHI3Z1(
.number_in1(VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1_number),
.read_add1(VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1_read_add),
.vmstubin(VMS_L5D3PHI3Z1n5_ME_L3L4_L5D3PHI3Z1),
.number_in2(VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1_number),
.read_add2(VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI3Z1_ME_L3L4_L5D3PHI3Z1),
.matchout(ME_L3L4_L5D3PHI3Z1_CM_L3L4_L5D3PHI3Z1),
.valid_data(ME_L3L4_L5D3PHI3Z1_CM_L3L4_L5D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D3PHI3Z2(
.number_in1(VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2_number),
.read_add1(VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2_read_add),
.vmstubin(VMS_L5D3PHI3Z2n5_ME_L3L4_L5D3PHI3Z2),
.number_in2(VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2_number),
.read_add2(VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI3Z2_ME_L3L4_L5D3PHI3Z2),
.matchout(ME_L3L4_L5D3PHI3Z2_CM_L3L4_L5D3PHI3Z2),
.valid_data(ME_L3L4_L5D3PHI3Z2_CM_L3L4_L5D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D4PHI1Z1(
.number_in1(VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1_number),
.read_add1(VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1_read_add),
.vmstubin(VMS_L5D4PHI1Z1n5_ME_L3L4_L5D4PHI1Z1),
.number_in2(VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1_number),
.read_add2(VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI1Z1_ME_L3L4_L5D4PHI1Z1),
.matchout(ME_L3L4_L5D4PHI1Z1_CM_L3L4_L5D4PHI1Z1),
.valid_data(ME_L3L4_L5D4PHI1Z1_CM_L3L4_L5D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D4PHI1Z2(
.number_in1(VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2_number),
.read_add1(VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2_read_add),
.vmstubin(VMS_L5D4PHI1Z2n3_ME_L3L4_L5D4PHI1Z2),
.number_in2(VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2_number),
.read_add2(VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI1Z2_ME_L3L4_L5D4PHI1Z2),
.matchout(ME_L3L4_L5D4PHI1Z2_CM_L3L4_L5D4PHI1Z2),
.valid_data(ME_L3L4_L5D4PHI1Z2_CM_L3L4_L5D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D4PHI2Z1(
.number_in1(VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1_number),
.read_add1(VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1_read_add),
.vmstubin(VMS_L5D4PHI2Z1n5_ME_L3L4_L5D4PHI2Z1),
.number_in2(VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1_number),
.read_add2(VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI2Z1_ME_L3L4_L5D4PHI2Z1),
.matchout(ME_L3L4_L5D4PHI2Z1_CM_L3L4_L5D4PHI2Z1),
.valid_data(ME_L3L4_L5D4PHI2Z1_CM_L3L4_L5D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D4PHI2Z2(
.number_in1(VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2_number),
.read_add1(VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2_read_add),
.vmstubin(VMS_L5D4PHI2Z2n3_ME_L3L4_L5D4PHI2Z2),
.number_in2(VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2_number),
.read_add2(VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI2Z2_ME_L3L4_L5D4PHI2Z2),
.matchout(ME_L3L4_L5D4PHI2Z2_CM_L3L4_L5D4PHI2Z2),
.valid_data(ME_L3L4_L5D4PHI2Z2_CM_L3L4_L5D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D4PHI3Z1(
.number_in1(VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1_number),
.read_add1(VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1_read_add),
.vmstubin(VMS_L5D4PHI3Z1n5_ME_L3L4_L5D4PHI3Z1),
.number_in2(VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1_number),
.read_add2(VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI3Z1_ME_L3L4_L5D4PHI3Z1),
.matchout(ME_L3L4_L5D4PHI3Z1_CM_L3L4_L5D4PHI3Z1),
.valid_data(ME_L3L4_L5D4PHI3Z1_CM_L3L4_L5D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L5D4PHI3Z2(
.number_in1(VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2_number),
.read_add1(VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2_read_add),
.vmstubin(VMS_L5D4PHI3Z2n3_ME_L3L4_L5D4PHI3Z2),
.number_in2(VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2_number),
.read_add2(VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI3Z2_ME_L3L4_L5D4PHI3Z2),
.matchout(ME_L3L4_L5D4PHI3Z2_CM_L3L4_L5D4PHI3Z2),
.valid_data(ME_L3L4_L5D4PHI3Z2_CM_L3L4_L5D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D3PHI1Z1(
.number_in1(VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1_number),
.read_add1(VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1_read_add),
.vmstubin(VMS_L6D3PHI1Z1n2_ME_L3L4_L6D3PHI1Z1),
.number_in2(VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1_number),
.read_add2(VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI1Z1_ME_L3L4_L6D3PHI1Z1),
.matchout(ME_L3L4_L6D3PHI1Z1_CM_L3L4_L6D3PHI1Z1),
.valid_data(ME_L3L4_L6D3PHI1Z1_CM_L3L4_L6D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D3PHI1Z2(
.number_in1(VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2_number),
.read_add1(VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2_read_add),
.vmstubin(VMS_L6D3PHI1Z2n3_ME_L3L4_L6D3PHI1Z2),
.number_in2(VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2_number),
.read_add2(VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI1Z2_ME_L3L4_L6D3PHI1Z2),
.matchout(ME_L3L4_L6D3PHI1Z2_CM_L3L4_L6D3PHI1Z2),
.valid_data(ME_L3L4_L6D3PHI1Z2_CM_L3L4_L6D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D3PHI2Z1(
.number_in1(VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1_number),
.read_add1(VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1_read_add),
.vmstubin(VMS_L6D3PHI2Z1n3_ME_L3L4_L6D3PHI2Z1),
.number_in2(VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1_number),
.read_add2(VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI2Z1_ME_L3L4_L6D3PHI2Z1),
.matchout(ME_L3L4_L6D3PHI2Z1_CM_L3L4_L6D3PHI2Z1),
.valid_data(ME_L3L4_L6D3PHI2Z1_CM_L3L4_L6D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D3PHI2Z2(
.number_in1(VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2_number),
.read_add1(VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2_read_add),
.vmstubin(VMS_L6D3PHI2Z2n5_ME_L3L4_L6D3PHI2Z2),
.number_in2(VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2_number),
.read_add2(VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI2Z2_ME_L3L4_L6D3PHI2Z2),
.matchout(ME_L3L4_L6D3PHI2Z2_CM_L3L4_L6D3PHI2Z2),
.valid_data(ME_L3L4_L6D3PHI2Z2_CM_L3L4_L6D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D3PHI3Z1(
.number_in1(VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1_number),
.read_add1(VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1_read_add),
.vmstubin(VMS_L6D3PHI3Z1n3_ME_L3L4_L6D3PHI3Z1),
.number_in2(VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1_number),
.read_add2(VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI3Z1_ME_L3L4_L6D3PHI3Z1),
.matchout(ME_L3L4_L6D3PHI3Z1_CM_L3L4_L6D3PHI3Z1),
.valid_data(ME_L3L4_L6D3PHI3Z1_CM_L3L4_L6D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D3PHI3Z2(
.number_in1(VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2_number),
.read_add1(VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2_read_add),
.vmstubin(VMS_L6D3PHI3Z2n5_ME_L3L4_L6D3PHI3Z2),
.number_in2(VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2_number),
.read_add2(VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI3Z2_ME_L3L4_L6D3PHI3Z2),
.matchout(ME_L3L4_L6D3PHI3Z2_CM_L3L4_L6D3PHI3Z2),
.valid_data(ME_L3L4_L6D3PHI3Z2_CM_L3L4_L6D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D3PHI4Z1(
.number_in1(VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1_number),
.read_add1(VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1_read_add),
.vmstubin(VMS_L6D3PHI4Z1n2_ME_L3L4_L6D3PHI4Z1),
.number_in2(VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1_number),
.read_add2(VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI4Z1_ME_L3L4_L6D3PHI4Z1),
.matchout(ME_L3L4_L6D3PHI4Z1_CM_L3L4_L6D3PHI4Z1),
.valid_data(ME_L3L4_L6D3PHI4Z1_CM_L3L4_L6D3PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D3PHI4Z2(
.number_in1(VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2_number),
.read_add1(VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2_read_add),
.vmstubin(VMS_L6D3PHI4Z2n3_ME_L3L4_L6D3PHI4Z2),
.number_in2(VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2_number),
.read_add2(VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI4Z2_ME_L3L4_L6D3PHI4Z2),
.matchout(ME_L3L4_L6D3PHI4Z2_CM_L3L4_L6D3PHI4Z2),
.valid_data(ME_L3L4_L6D3PHI4Z2_CM_L3L4_L6D3PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D4PHI1Z1(
.number_in1(VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1_number),
.read_add1(VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1_read_add),
.vmstubin(VMS_L6D4PHI1Z1n3_ME_L3L4_L6D4PHI1Z1),
.number_in2(VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1_number),
.read_add2(VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI1Z1_ME_L3L4_L6D4PHI1Z1),
.matchout(ME_L3L4_L6D4PHI1Z1_CM_L3L4_L6D4PHI1Z1),
.valid_data(ME_L3L4_L6D4PHI1Z1_CM_L3L4_L6D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D4PHI1Z2(
.number_in1(VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2_number),
.read_add1(VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2_read_add),
.vmstubin(VMS_L6D4PHI1Z2n3_ME_L3L4_L6D4PHI1Z2),
.number_in2(VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2_number),
.read_add2(VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI1Z2_ME_L3L4_L6D4PHI1Z2),
.matchout(ME_L3L4_L6D4PHI1Z2_CM_L3L4_L6D4PHI1Z2),
.valid_data(ME_L3L4_L6D4PHI1Z2_CM_L3L4_L6D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D4PHI2Z1(
.number_in1(VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1_number),
.read_add1(VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1_read_add),
.vmstubin(VMS_L6D4PHI2Z1n5_ME_L3L4_L6D4PHI2Z1),
.number_in2(VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1_number),
.read_add2(VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI2Z1_ME_L3L4_L6D4PHI2Z1),
.matchout(ME_L3L4_L6D4PHI2Z1_CM_L3L4_L6D4PHI2Z1),
.valid_data(ME_L3L4_L6D4PHI2Z1_CM_L3L4_L6D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D4PHI2Z2(
.number_in1(VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2_number),
.read_add1(VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2_read_add),
.vmstubin(VMS_L6D4PHI2Z2n5_ME_L3L4_L6D4PHI2Z2),
.number_in2(VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2_number),
.read_add2(VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI2Z2_ME_L3L4_L6D4PHI2Z2),
.matchout(ME_L3L4_L6D4PHI2Z2_CM_L3L4_L6D4PHI2Z2),
.valid_data(ME_L3L4_L6D4PHI2Z2_CM_L3L4_L6D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D4PHI3Z1(
.number_in1(VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1_number),
.read_add1(VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1_read_add),
.vmstubin(VMS_L6D4PHI3Z1n5_ME_L3L4_L6D4PHI3Z1),
.number_in2(VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1_number),
.read_add2(VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI3Z1_ME_L3L4_L6D4PHI3Z1),
.matchout(ME_L3L4_L6D4PHI3Z1_CM_L3L4_L6D4PHI3Z1),
.valid_data(ME_L3L4_L6D4PHI3Z1_CM_L3L4_L6D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D4PHI3Z2(
.number_in1(VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2_number),
.read_add1(VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2_read_add),
.vmstubin(VMS_L6D4PHI3Z2n5_ME_L3L4_L6D4PHI3Z2),
.number_in2(VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2_number),
.read_add2(VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI3Z2_ME_L3L4_L6D4PHI3Z2),
.matchout(ME_L3L4_L6D4PHI3Z2_CM_L3L4_L6D4PHI3Z2),
.valid_data(ME_L3L4_L6D4PHI3Z2_CM_L3L4_L6D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D4PHI4Z1(
.number_in1(VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1_number),
.read_add1(VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1_read_add),
.vmstubin(VMS_L6D4PHI4Z1n3_ME_L3L4_L6D4PHI4Z1),
.number_in2(VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1_number),
.read_add2(VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI4Z1_ME_L3L4_L6D4PHI4Z1),
.matchout(ME_L3L4_L6D4PHI4Z1_CM_L3L4_L6D4PHI4Z1),
.valid_data(ME_L3L4_L6D4PHI4Z1_CM_L3L4_L6D4PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L3L4_L6D4PHI4Z2(
.number_in1(VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2_number),
.read_add1(VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2_read_add),
.vmstubin(VMS_L6D4PHI4Z2n3_ME_L3L4_L6D4PHI4Z2),
.number_in2(VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2_number),
.read_add2(VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI4Z2_ME_L3L4_L6D4PHI4Z2),
.matchout(ME_L3L4_L6D4PHI4Z2_CM_L3L4_L6D4PHI4Z2),
.valid_data(ME_L3L4_L6D4PHI4Z2_CM_L3L4_L6D4PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D3PHI1Z1(
.number_in1(VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1_number),
.read_add1(VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1_read_add),
.vmstubin(VMS_L3D3PHI1Z1n5_ME_L1L2_L3D3PHI1Z1),
.number_in2(VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1_number),
.read_add2(VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI1Z1_ME_L1L2_L3D3PHI1Z1),
.matchout(ME_L1L2_L3D3PHI1Z1_CM_L1L2_L3D3PHI1Z1),
.valid_data(ME_L1L2_L3D3PHI1Z1_CM_L1L2_L3D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D3PHI1Z2(
.number_in1(VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2_number),
.read_add1(VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2_read_add),
.vmstubin(VMS_L3D3PHI1Z2n5_ME_L1L2_L3D3PHI1Z2),
.number_in2(VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2_number),
.read_add2(VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI1Z2_ME_L1L2_L3D3PHI1Z2),
.matchout(ME_L1L2_L3D3PHI1Z2_CM_L1L2_L3D3PHI1Z2),
.valid_data(ME_L1L2_L3D3PHI1Z2_CM_L1L2_L3D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D3PHI2Z1(
.number_in1(VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1_number),
.read_add1(VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1_read_add),
.vmstubin(VMS_L3D3PHI2Z1n5_ME_L1L2_L3D3PHI2Z1),
.number_in2(VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1_number),
.read_add2(VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI2Z1_ME_L1L2_L3D3PHI2Z1),
.matchout(ME_L1L2_L3D3PHI2Z1_CM_L1L2_L3D3PHI2Z1),
.valid_data(ME_L1L2_L3D3PHI2Z1_CM_L1L2_L3D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D3PHI2Z2(
.number_in1(VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2_number),
.read_add1(VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2_read_add),
.vmstubin(VMS_L3D3PHI2Z2n5_ME_L1L2_L3D3PHI2Z2),
.number_in2(VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2_number),
.read_add2(VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI2Z2_ME_L1L2_L3D3PHI2Z2),
.matchout(ME_L1L2_L3D3PHI2Z2_CM_L1L2_L3D3PHI2Z2),
.valid_data(ME_L1L2_L3D3PHI2Z2_CM_L1L2_L3D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D3PHI3Z1(
.number_in1(VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1_number),
.read_add1(VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1_read_add),
.vmstubin(VMS_L3D3PHI3Z1n5_ME_L1L2_L3D3PHI3Z1),
.number_in2(VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1_number),
.read_add2(VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI3Z1_ME_L1L2_L3D3PHI3Z1),
.matchout(ME_L1L2_L3D3PHI3Z1_CM_L1L2_L3D3PHI3Z1),
.valid_data(ME_L1L2_L3D3PHI3Z1_CM_L1L2_L3D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D3PHI3Z2(
.number_in1(VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2_number),
.read_add1(VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2_read_add),
.vmstubin(VMS_L3D3PHI3Z2n5_ME_L1L2_L3D3PHI3Z2),
.number_in2(VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2_number),
.read_add2(VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI3Z2_ME_L1L2_L3D3PHI3Z2),
.matchout(ME_L1L2_L3D3PHI3Z2_CM_L1L2_L3D3PHI3Z2),
.valid_data(ME_L1L2_L3D3PHI3Z2_CM_L1L2_L3D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D4PHI1Z1(
.number_in1(VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1_number),
.read_add1(VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1_read_add),
.vmstubin(VMS_L3D4PHI1Z1n5_ME_L1L2_L3D4PHI1Z1),
.number_in2(VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1_number),
.read_add2(VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI1Z1_ME_L1L2_L3D4PHI1Z1),
.matchout(ME_L1L2_L3D4PHI1Z1_CM_L1L2_L3D4PHI1Z1),
.valid_data(ME_L1L2_L3D4PHI1Z1_CM_L1L2_L3D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D4PHI1Z2(
.number_in1(VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2_number),
.read_add1(VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2_read_add),
.vmstubin(VMS_L3D4PHI1Z2n3_ME_L1L2_L3D4PHI1Z2),
.number_in2(VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2_number),
.read_add2(VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI1Z2_ME_L1L2_L3D4PHI1Z2),
.matchout(ME_L1L2_L3D4PHI1Z2_CM_L1L2_L3D4PHI1Z2),
.valid_data(ME_L1L2_L3D4PHI1Z2_CM_L1L2_L3D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D4PHI2Z1(
.number_in1(VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1_number),
.read_add1(VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1_read_add),
.vmstubin(VMS_L3D4PHI2Z1n5_ME_L1L2_L3D4PHI2Z1),
.number_in2(VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1_number),
.read_add2(VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI2Z1_ME_L1L2_L3D4PHI2Z1),
.matchout(ME_L1L2_L3D4PHI2Z1_CM_L1L2_L3D4PHI2Z1),
.valid_data(ME_L1L2_L3D4PHI2Z1_CM_L1L2_L3D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D4PHI2Z2(
.number_in1(VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2_number),
.read_add1(VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2_read_add),
.vmstubin(VMS_L3D4PHI2Z2n3_ME_L1L2_L3D4PHI2Z2),
.number_in2(VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2_number),
.read_add2(VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI2Z2_ME_L1L2_L3D4PHI2Z2),
.matchout(ME_L1L2_L3D4PHI2Z2_CM_L1L2_L3D4PHI2Z2),
.valid_data(ME_L1L2_L3D4PHI2Z2_CM_L1L2_L3D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D4PHI3Z1(
.number_in1(VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1_number),
.read_add1(VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1_read_add),
.vmstubin(VMS_L3D4PHI3Z1n5_ME_L1L2_L3D4PHI3Z1),
.number_in2(VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1_number),
.read_add2(VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI3Z1_ME_L1L2_L3D4PHI3Z1),
.matchout(ME_L1L2_L3D4PHI3Z1_CM_L1L2_L3D4PHI3Z1),
.valid_data(ME_L1L2_L3D4PHI3Z1_CM_L1L2_L3D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L3D4PHI3Z2(
.number_in1(VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2_number),
.read_add1(VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2_read_add),
.vmstubin(VMS_L3D4PHI3Z2n3_ME_L1L2_L3D4PHI3Z2),
.number_in2(VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2_number),
.read_add2(VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI3Z2_ME_L1L2_L3D4PHI3Z2),
.matchout(ME_L1L2_L3D4PHI3Z2_CM_L1L2_L3D4PHI3Z2),
.valid_data(ME_L1L2_L3D4PHI3Z2_CM_L1L2_L3D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D3PHI1Z1(
.number_in1(VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1_number),
.read_add1(VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1_read_add),
.vmstubin(VMS_L4D3PHI1Z1n2_ME_L1L2_L4D3PHI1Z1),
.number_in2(VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1_number),
.read_add2(VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI1Z1_ME_L1L2_L4D3PHI1Z1),
.matchout(ME_L1L2_L4D3PHI1Z1_CM_L1L2_L4D3PHI1Z1),
.valid_data(ME_L1L2_L4D3PHI1Z1_CM_L1L2_L4D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D3PHI1Z2(
.number_in1(VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2_number),
.read_add1(VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2_read_add),
.vmstubin(VMS_L4D3PHI1Z2n3_ME_L1L2_L4D3PHI1Z2),
.number_in2(VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2_number),
.read_add2(VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI1Z2_ME_L1L2_L4D3PHI1Z2),
.matchout(ME_L1L2_L4D3PHI1Z2_CM_L1L2_L4D3PHI1Z2),
.valid_data(ME_L1L2_L4D3PHI1Z2_CM_L1L2_L4D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D3PHI2Z1(
.number_in1(VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1_number),
.read_add1(VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1_read_add),
.vmstubin(VMS_L4D3PHI2Z1n3_ME_L1L2_L4D3PHI2Z1),
.number_in2(VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1_number),
.read_add2(VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI2Z1_ME_L1L2_L4D3PHI2Z1),
.matchout(ME_L1L2_L4D3PHI2Z1_CM_L1L2_L4D3PHI2Z1),
.valid_data(ME_L1L2_L4D3PHI2Z1_CM_L1L2_L4D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D3PHI2Z2(
.number_in1(VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2_number),
.read_add1(VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2_read_add),
.vmstubin(VMS_L4D3PHI2Z2n5_ME_L1L2_L4D3PHI2Z2),
.number_in2(VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2_number),
.read_add2(VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI2Z2_ME_L1L2_L4D3PHI2Z2),
.matchout(ME_L1L2_L4D3PHI2Z2_CM_L1L2_L4D3PHI2Z2),
.valid_data(ME_L1L2_L4D3PHI2Z2_CM_L1L2_L4D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D3PHI3Z1(
.number_in1(VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1_number),
.read_add1(VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1_read_add),
.vmstubin(VMS_L4D3PHI3Z1n3_ME_L1L2_L4D3PHI3Z1),
.number_in2(VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1_number),
.read_add2(VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI3Z1_ME_L1L2_L4D3PHI3Z1),
.matchout(ME_L1L2_L4D3PHI3Z1_CM_L1L2_L4D3PHI3Z1),
.valid_data(ME_L1L2_L4D3PHI3Z1_CM_L1L2_L4D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D3PHI3Z2(
.number_in1(VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2_number),
.read_add1(VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2_read_add),
.vmstubin(VMS_L4D3PHI3Z2n5_ME_L1L2_L4D3PHI3Z2),
.number_in2(VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2_number),
.read_add2(VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI3Z2_ME_L1L2_L4D3PHI3Z2),
.matchout(ME_L1L2_L4D3PHI3Z2_CM_L1L2_L4D3PHI3Z2),
.valid_data(ME_L1L2_L4D3PHI3Z2_CM_L1L2_L4D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D3PHI4Z1(
.number_in1(VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1_number),
.read_add1(VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1_read_add),
.vmstubin(VMS_L4D3PHI4Z1n2_ME_L1L2_L4D3PHI4Z1),
.number_in2(VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1_number),
.read_add2(VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI4Z1_ME_L1L2_L4D3PHI4Z1),
.matchout(ME_L1L2_L4D3PHI4Z1_CM_L1L2_L4D3PHI4Z1),
.valid_data(ME_L1L2_L4D3PHI4Z1_CM_L1L2_L4D3PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D3PHI4Z2(
.number_in1(VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2_number),
.read_add1(VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2_read_add),
.vmstubin(VMS_L4D3PHI4Z2n3_ME_L1L2_L4D3PHI4Z2),
.number_in2(VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2_number),
.read_add2(VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI4Z2_ME_L1L2_L4D3PHI4Z2),
.matchout(ME_L1L2_L4D3PHI4Z2_CM_L1L2_L4D3PHI4Z2),
.valid_data(ME_L1L2_L4D3PHI4Z2_CM_L1L2_L4D3PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D4PHI1Z1(
.number_in1(VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1_number),
.read_add1(VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1_read_add),
.vmstubin(VMS_L4D4PHI1Z1n3_ME_L1L2_L4D4PHI1Z1),
.number_in2(VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1_number),
.read_add2(VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI1Z1_ME_L1L2_L4D4PHI1Z1),
.matchout(ME_L1L2_L4D4PHI1Z1_CM_L1L2_L4D4PHI1Z1),
.valid_data(ME_L1L2_L4D4PHI1Z1_CM_L1L2_L4D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D4PHI1Z2(
.number_in1(VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2_number),
.read_add1(VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2_read_add),
.vmstubin(VMS_L4D4PHI1Z2n3_ME_L1L2_L4D4PHI1Z2),
.number_in2(VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2_number),
.read_add2(VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI1Z2_ME_L1L2_L4D4PHI1Z2),
.matchout(ME_L1L2_L4D4PHI1Z2_CM_L1L2_L4D4PHI1Z2),
.valid_data(ME_L1L2_L4D4PHI1Z2_CM_L1L2_L4D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D4PHI2Z1(
.number_in1(VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1_number),
.read_add1(VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1_read_add),
.vmstubin(VMS_L4D4PHI2Z1n5_ME_L1L2_L4D4PHI2Z1),
.number_in2(VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1_number),
.read_add2(VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI2Z1_ME_L1L2_L4D4PHI2Z1),
.matchout(ME_L1L2_L4D4PHI2Z1_CM_L1L2_L4D4PHI2Z1),
.valid_data(ME_L1L2_L4D4PHI2Z1_CM_L1L2_L4D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D4PHI2Z2(
.number_in1(VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2_number),
.read_add1(VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2_read_add),
.vmstubin(VMS_L4D4PHI2Z2n5_ME_L1L2_L4D4PHI2Z2),
.number_in2(VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2_number),
.read_add2(VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI2Z2_ME_L1L2_L4D4PHI2Z2),
.matchout(ME_L1L2_L4D4PHI2Z2_CM_L1L2_L4D4PHI2Z2),
.valid_data(ME_L1L2_L4D4PHI2Z2_CM_L1L2_L4D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D4PHI3Z1(
.number_in1(VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1_number),
.read_add1(VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1_read_add),
.vmstubin(VMS_L4D4PHI3Z1n5_ME_L1L2_L4D4PHI3Z1),
.number_in2(VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1_number),
.read_add2(VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI3Z1_ME_L1L2_L4D4PHI3Z1),
.matchout(ME_L1L2_L4D4PHI3Z1_CM_L1L2_L4D4PHI3Z1),
.valid_data(ME_L1L2_L4D4PHI3Z1_CM_L1L2_L4D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D4PHI3Z2(
.number_in1(VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2_number),
.read_add1(VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2_read_add),
.vmstubin(VMS_L4D4PHI3Z2n5_ME_L1L2_L4D4PHI3Z2),
.number_in2(VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2_number),
.read_add2(VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI3Z2_ME_L1L2_L4D4PHI3Z2),
.matchout(ME_L1L2_L4D4PHI3Z2_CM_L1L2_L4D4PHI3Z2),
.valid_data(ME_L1L2_L4D4PHI3Z2_CM_L1L2_L4D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D4PHI4Z1(
.number_in1(VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1_number),
.read_add1(VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1_read_add),
.vmstubin(VMS_L4D4PHI4Z1n3_ME_L1L2_L4D4PHI4Z1),
.number_in2(VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1_number),
.read_add2(VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI4Z1_ME_L1L2_L4D4PHI4Z1),
.matchout(ME_L1L2_L4D4PHI4Z1_CM_L1L2_L4D4PHI4Z1),
.valid_data(ME_L1L2_L4D4PHI4Z1_CM_L1L2_L4D4PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L4D4PHI4Z2(
.number_in1(VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2_number),
.read_add1(VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2_read_add),
.vmstubin(VMS_L4D4PHI4Z2n3_ME_L1L2_L4D4PHI4Z2),
.number_in2(VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2_number),
.read_add2(VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI4Z2_ME_L1L2_L4D4PHI4Z2),
.matchout(ME_L1L2_L4D4PHI4Z2_CM_L1L2_L4D4PHI4Z2),
.valid_data(ME_L1L2_L4D4PHI4Z2_CM_L1L2_L4D4PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D3PHI1Z1(
.number_in1(VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1_number),
.read_add1(VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1_read_add),
.vmstubin(VMS_L5D3PHI1Z1n6_ME_L1L2_L5D3PHI1Z1),
.number_in2(VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1_number),
.read_add2(VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI1Z1_ME_L1L2_L5D3PHI1Z1),
.matchout(ME_L1L2_L5D3PHI1Z1_CM_L1L2_L5D3PHI1Z1),
.valid_data(ME_L1L2_L5D3PHI1Z1_CM_L1L2_L5D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D3PHI1Z2(
.number_in1(VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2_number),
.read_add1(VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2_read_add),
.vmstubin(VMS_L5D3PHI1Z2n6_ME_L1L2_L5D3PHI1Z2),
.number_in2(VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2_number),
.read_add2(VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI1Z2_ME_L1L2_L5D3PHI1Z2),
.matchout(ME_L1L2_L5D3PHI1Z2_CM_L1L2_L5D3PHI1Z2),
.valid_data(ME_L1L2_L5D3PHI1Z2_CM_L1L2_L5D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D3PHI2Z1(
.number_in1(VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1_number),
.read_add1(VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1_read_add),
.vmstubin(VMS_L5D3PHI2Z1n6_ME_L1L2_L5D3PHI2Z1),
.number_in2(VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1_number),
.read_add2(VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI2Z1_ME_L1L2_L5D3PHI2Z1),
.matchout(ME_L1L2_L5D3PHI2Z1_CM_L1L2_L5D3PHI2Z1),
.valid_data(ME_L1L2_L5D3PHI2Z1_CM_L1L2_L5D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D3PHI2Z2(
.number_in1(VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2_number),
.read_add1(VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2_read_add),
.vmstubin(VMS_L5D3PHI2Z2n6_ME_L1L2_L5D3PHI2Z2),
.number_in2(VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2_number),
.read_add2(VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI2Z2_ME_L1L2_L5D3PHI2Z2),
.matchout(ME_L1L2_L5D3PHI2Z2_CM_L1L2_L5D3PHI2Z2),
.valid_data(ME_L1L2_L5D3PHI2Z2_CM_L1L2_L5D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D3PHI3Z1(
.number_in1(VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1_number),
.read_add1(VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1_read_add),
.vmstubin(VMS_L5D3PHI3Z1n6_ME_L1L2_L5D3PHI3Z1),
.number_in2(VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1_number),
.read_add2(VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI3Z1_ME_L1L2_L5D3PHI3Z1),
.matchout(ME_L1L2_L5D3PHI3Z1_CM_L1L2_L5D3PHI3Z1),
.valid_data(ME_L1L2_L5D3PHI3Z1_CM_L1L2_L5D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D3PHI3Z2(
.number_in1(VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2_number),
.read_add1(VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2_read_add),
.vmstubin(VMS_L5D3PHI3Z2n6_ME_L1L2_L5D3PHI3Z2),
.number_in2(VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2_number),
.read_add2(VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI3Z2_ME_L1L2_L5D3PHI3Z2),
.matchout(ME_L1L2_L5D3PHI3Z2_CM_L1L2_L5D3PHI3Z2),
.valid_data(ME_L1L2_L5D3PHI3Z2_CM_L1L2_L5D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D4PHI1Z1(
.number_in1(VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1_number),
.read_add1(VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1_read_add),
.vmstubin(VMS_L5D4PHI1Z1n6_ME_L1L2_L5D4PHI1Z1),
.number_in2(VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1_number),
.read_add2(VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI1Z1_ME_L1L2_L5D4PHI1Z1),
.matchout(ME_L1L2_L5D4PHI1Z1_CM_L1L2_L5D4PHI1Z1),
.valid_data(ME_L1L2_L5D4PHI1Z1_CM_L1L2_L5D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D4PHI1Z2(
.number_in1(VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2_number),
.read_add1(VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2_read_add),
.vmstubin(VMS_L5D4PHI1Z2n4_ME_L1L2_L5D4PHI1Z2),
.number_in2(VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2_number),
.read_add2(VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI1Z2_ME_L1L2_L5D4PHI1Z2),
.matchout(ME_L1L2_L5D4PHI1Z2_CM_L1L2_L5D4PHI1Z2),
.valid_data(ME_L1L2_L5D4PHI1Z2_CM_L1L2_L5D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D4PHI2Z1(
.number_in1(VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1_number),
.read_add1(VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1_read_add),
.vmstubin(VMS_L5D4PHI2Z1n6_ME_L1L2_L5D4PHI2Z1),
.number_in2(VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1_number),
.read_add2(VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI2Z1_ME_L1L2_L5D4PHI2Z1),
.matchout(ME_L1L2_L5D4PHI2Z1_CM_L1L2_L5D4PHI2Z1),
.valid_data(ME_L1L2_L5D4PHI2Z1_CM_L1L2_L5D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D4PHI2Z2(
.number_in1(VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2_number),
.read_add1(VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2_read_add),
.vmstubin(VMS_L5D4PHI2Z2n4_ME_L1L2_L5D4PHI2Z2),
.number_in2(VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2_number),
.read_add2(VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI2Z2_ME_L1L2_L5D4PHI2Z2),
.matchout(ME_L1L2_L5D4PHI2Z2_CM_L1L2_L5D4PHI2Z2),
.valid_data(ME_L1L2_L5D4PHI2Z2_CM_L1L2_L5D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D4PHI3Z1(
.number_in1(VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1_number),
.read_add1(VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1_read_add),
.vmstubin(VMS_L5D4PHI3Z1n6_ME_L1L2_L5D4PHI3Z1),
.number_in2(VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1_number),
.read_add2(VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI3Z1_ME_L1L2_L5D4PHI3Z1),
.matchout(ME_L1L2_L5D4PHI3Z1_CM_L1L2_L5D4PHI3Z1),
.valid_data(ME_L1L2_L5D4PHI3Z1_CM_L1L2_L5D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L5D4PHI3Z2(
.number_in1(VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2_number),
.read_add1(VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2_read_add),
.vmstubin(VMS_L5D4PHI3Z2n4_ME_L1L2_L5D4PHI3Z2),
.number_in2(VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2_number),
.read_add2(VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI3Z2_ME_L1L2_L5D4PHI3Z2),
.matchout(ME_L1L2_L5D4PHI3Z2_CM_L1L2_L5D4PHI3Z2),
.valid_data(ME_L1L2_L5D4PHI3Z2_CM_L1L2_L5D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D3PHI1Z1(
.number_in1(VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1_number),
.read_add1(VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1_read_add),
.vmstubin(VMS_L6D3PHI1Z1n3_ME_L1L2_L6D3PHI1Z1),
.number_in2(VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1_number),
.read_add2(VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI1Z1_ME_L1L2_L6D3PHI1Z1),
.matchout(ME_L1L2_L6D3PHI1Z1_CM_L1L2_L6D3PHI1Z1),
.valid_data(ME_L1L2_L6D3PHI1Z1_CM_L1L2_L6D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D3PHI1Z2(
.number_in1(VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2_number),
.read_add1(VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2_read_add),
.vmstubin(VMS_L6D3PHI1Z2n4_ME_L1L2_L6D3PHI1Z2),
.number_in2(VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2_number),
.read_add2(VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI1Z2_ME_L1L2_L6D3PHI1Z2),
.matchout(ME_L1L2_L6D3PHI1Z2_CM_L1L2_L6D3PHI1Z2),
.valid_data(ME_L1L2_L6D3PHI1Z2_CM_L1L2_L6D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D3PHI2Z1(
.number_in1(VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1_number),
.read_add1(VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1_read_add),
.vmstubin(VMS_L6D3PHI2Z1n4_ME_L1L2_L6D3PHI2Z1),
.number_in2(VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1_number),
.read_add2(VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI2Z1_ME_L1L2_L6D3PHI2Z1),
.matchout(ME_L1L2_L6D3PHI2Z1_CM_L1L2_L6D3PHI2Z1),
.valid_data(ME_L1L2_L6D3PHI2Z1_CM_L1L2_L6D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D3PHI2Z2(
.number_in1(VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2_number),
.read_add1(VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2_read_add),
.vmstubin(VMS_L6D3PHI2Z2n6_ME_L1L2_L6D3PHI2Z2),
.number_in2(VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2_number),
.read_add2(VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI2Z2_ME_L1L2_L6D3PHI2Z2),
.matchout(ME_L1L2_L6D3PHI2Z2_CM_L1L2_L6D3PHI2Z2),
.valid_data(ME_L1L2_L6D3PHI2Z2_CM_L1L2_L6D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D3PHI3Z1(
.number_in1(VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1_number),
.read_add1(VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1_read_add),
.vmstubin(VMS_L6D3PHI3Z1n4_ME_L1L2_L6D3PHI3Z1),
.number_in2(VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1_number),
.read_add2(VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI3Z1_ME_L1L2_L6D3PHI3Z1),
.matchout(ME_L1L2_L6D3PHI3Z1_CM_L1L2_L6D3PHI3Z1),
.valid_data(ME_L1L2_L6D3PHI3Z1_CM_L1L2_L6D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D3PHI3Z2(
.number_in1(VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2_number),
.read_add1(VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2_read_add),
.vmstubin(VMS_L6D3PHI3Z2n6_ME_L1L2_L6D3PHI3Z2),
.number_in2(VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2_number),
.read_add2(VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI3Z2_ME_L1L2_L6D3PHI3Z2),
.matchout(ME_L1L2_L6D3PHI3Z2_CM_L1L2_L6D3PHI3Z2),
.valid_data(ME_L1L2_L6D3PHI3Z2_CM_L1L2_L6D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D3PHI4Z1(
.number_in1(VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1_number),
.read_add1(VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1_read_add),
.vmstubin(VMS_L6D3PHI4Z1n3_ME_L1L2_L6D3PHI4Z1),
.number_in2(VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1_number),
.read_add2(VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI4Z1_ME_L1L2_L6D3PHI4Z1),
.matchout(ME_L1L2_L6D3PHI4Z1_CM_L1L2_L6D3PHI4Z1),
.valid_data(ME_L1L2_L6D3PHI4Z1_CM_L1L2_L6D3PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D3PHI4Z2(
.number_in1(VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2_number),
.read_add1(VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2_read_add),
.vmstubin(VMS_L6D3PHI4Z2n4_ME_L1L2_L6D3PHI4Z2),
.number_in2(VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2_number),
.read_add2(VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI4Z2_ME_L1L2_L6D3PHI4Z2),
.matchout(ME_L1L2_L6D3PHI4Z2_CM_L1L2_L6D3PHI4Z2),
.valid_data(ME_L1L2_L6D3PHI4Z2_CM_L1L2_L6D3PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D4PHI1Z1(
.number_in1(VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1_number),
.read_add1(VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1_read_add),
.vmstubin(VMS_L6D4PHI1Z1n4_ME_L1L2_L6D4PHI1Z1),
.number_in2(VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1_number),
.read_add2(VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI1Z1_ME_L1L2_L6D4PHI1Z1),
.matchout(ME_L1L2_L6D4PHI1Z1_CM_L1L2_L6D4PHI1Z1),
.valid_data(ME_L1L2_L6D4PHI1Z1_CM_L1L2_L6D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D4PHI1Z2(
.number_in1(VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2_number),
.read_add1(VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2_read_add),
.vmstubin(VMS_L6D4PHI1Z2n4_ME_L1L2_L6D4PHI1Z2),
.number_in2(VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2_number),
.read_add2(VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI1Z2_ME_L1L2_L6D4PHI1Z2),
.matchout(ME_L1L2_L6D4PHI1Z2_CM_L1L2_L6D4PHI1Z2),
.valid_data(ME_L1L2_L6D4PHI1Z2_CM_L1L2_L6D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D4PHI2Z1(
.number_in1(VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1_number),
.read_add1(VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1_read_add),
.vmstubin(VMS_L6D4PHI2Z1n6_ME_L1L2_L6D4PHI2Z1),
.number_in2(VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1_number),
.read_add2(VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI2Z1_ME_L1L2_L6D4PHI2Z1),
.matchout(ME_L1L2_L6D4PHI2Z1_CM_L1L2_L6D4PHI2Z1),
.valid_data(ME_L1L2_L6D4PHI2Z1_CM_L1L2_L6D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D4PHI2Z2(
.number_in1(VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2_number),
.read_add1(VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2_read_add),
.vmstubin(VMS_L6D4PHI2Z2n6_ME_L1L2_L6D4PHI2Z2),
.number_in2(VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2_number),
.read_add2(VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI2Z2_ME_L1L2_L6D4PHI2Z2),
.matchout(ME_L1L2_L6D4PHI2Z2_CM_L1L2_L6D4PHI2Z2),
.valid_data(ME_L1L2_L6D4PHI2Z2_CM_L1L2_L6D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D4PHI3Z1(
.number_in1(VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1_number),
.read_add1(VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1_read_add),
.vmstubin(VMS_L6D4PHI3Z1n6_ME_L1L2_L6D4PHI3Z1),
.number_in2(VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1_number),
.read_add2(VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI3Z1_ME_L1L2_L6D4PHI3Z1),
.matchout(ME_L1L2_L6D4PHI3Z1_CM_L1L2_L6D4PHI3Z1),
.valid_data(ME_L1L2_L6D4PHI3Z1_CM_L1L2_L6D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D4PHI3Z2(
.number_in1(VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2_number),
.read_add1(VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2_read_add),
.vmstubin(VMS_L6D4PHI3Z2n6_ME_L1L2_L6D4PHI3Z2),
.number_in2(VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2_number),
.read_add2(VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI3Z2_ME_L1L2_L6D4PHI3Z2),
.matchout(ME_L1L2_L6D4PHI3Z2_CM_L1L2_L6D4PHI3Z2),
.valid_data(ME_L1L2_L6D4PHI3Z2_CM_L1L2_L6D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D4PHI4Z1(
.number_in1(VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1_number),
.read_add1(VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1_read_add),
.vmstubin(VMS_L6D4PHI4Z1n4_ME_L1L2_L6D4PHI4Z1),
.number_in2(VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1_number),
.read_add2(VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI4Z1_ME_L1L2_L6D4PHI4Z1),
.matchout(ME_L1L2_L6D4PHI4Z1_CM_L1L2_L6D4PHI4Z1),
.valid_data(ME_L1L2_L6D4PHI4Z1_CM_L1L2_L6D4PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L1L2_L6D4PHI4Z2(
.number_in1(VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2_number),
.read_add1(VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2_read_add),
.vmstubin(VMS_L6D4PHI4Z2n4_ME_L1L2_L6D4PHI4Z2),
.number_in2(VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2_number),
.read_add2(VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI4Z2_ME_L1L2_L6D4PHI4Z2),
.matchout(ME_L1L2_L6D4PHI4Z2_CM_L1L2_L6D4PHI4Z2),
.valid_data(ME_L1L2_L6D4PHI4Z2_CM_L1L2_L6D4PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D3PHI1Z1(
.number_in1(VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1_number),
.read_add1(VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1_read_add),
.vmstubin(VMS_L1D3PHI1Z1n8_ME_L5L6_L1D3PHI1Z1),
.number_in2(VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1_number),
.read_add2(VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI1Z1_ME_L5L6_L1D3PHI1Z1),
.matchout(ME_L5L6_L1D3PHI1Z1_CM_L5L6_L1D3PHI1Z1),
.valid_data(ME_L5L6_L1D3PHI1Z1_CM_L5L6_L1D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D3PHI1Z2(
.number_in1(VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2_number),
.read_add1(VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2_read_add),
.vmstubin(VMS_L1D3PHI1Z2n8_ME_L5L6_L1D3PHI1Z2),
.number_in2(VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2_number),
.read_add2(VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI1Z2_ME_L5L6_L1D3PHI1Z2),
.matchout(ME_L5L6_L1D3PHI1Z2_CM_L5L6_L1D3PHI1Z2),
.valid_data(ME_L5L6_L1D3PHI1Z2_CM_L5L6_L1D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D3PHI2Z1(
.number_in1(VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1_number),
.read_add1(VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1_read_add),
.vmstubin(VMS_L1D3PHI2Z1n8_ME_L5L6_L1D3PHI2Z1),
.number_in2(VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1_number),
.read_add2(VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI2Z1_ME_L5L6_L1D3PHI2Z1),
.matchout(ME_L5L6_L1D3PHI2Z1_CM_L5L6_L1D3PHI2Z1),
.valid_data(ME_L5L6_L1D3PHI2Z1_CM_L5L6_L1D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D3PHI2Z2(
.number_in1(VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2_number),
.read_add1(VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2_read_add),
.vmstubin(VMS_L1D3PHI2Z2n8_ME_L5L6_L1D3PHI2Z2),
.number_in2(VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2_number),
.read_add2(VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI2Z2_ME_L5L6_L1D3PHI2Z2),
.matchout(ME_L5L6_L1D3PHI2Z2_CM_L5L6_L1D3PHI2Z2),
.valid_data(ME_L5L6_L1D3PHI2Z2_CM_L5L6_L1D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D3PHI3Z1(
.number_in1(VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1_number),
.read_add1(VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1_read_add),
.vmstubin(VMS_L1D3PHI3Z1n8_ME_L5L6_L1D3PHI3Z1),
.number_in2(VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1_number),
.read_add2(VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI3Z1_ME_L5L6_L1D3PHI3Z1),
.matchout(ME_L5L6_L1D3PHI3Z1_CM_L5L6_L1D3PHI3Z1),
.valid_data(ME_L5L6_L1D3PHI3Z1_CM_L5L6_L1D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D3PHI3Z2(
.number_in1(VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2_number),
.read_add1(VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2_read_add),
.vmstubin(VMS_L1D3PHI3Z2n8_ME_L5L6_L1D3PHI3Z2),
.number_in2(VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2_number),
.read_add2(VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI3Z2_ME_L5L6_L1D3PHI3Z2),
.matchout(ME_L5L6_L1D3PHI3Z2_CM_L5L6_L1D3PHI3Z2),
.valid_data(ME_L5L6_L1D3PHI3Z2_CM_L5L6_L1D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D4PHI1Z1(
.number_in1(VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1_number),
.read_add1(VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1_read_add),
.vmstubin(VMS_L1D4PHI1Z1n4_ME_L5L6_L1D4PHI1Z1),
.number_in2(VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1_number),
.read_add2(VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI1Z1_ME_L5L6_L1D4PHI1Z1),
.matchout(ME_L5L6_L1D4PHI1Z1_CM_L5L6_L1D4PHI1Z1),
.valid_data(ME_L5L6_L1D4PHI1Z1_CM_L5L6_L1D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D4PHI1Z2(
.number_in1(VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2_number),
.read_add1(VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2_read_add),
.vmstubin(VMS_L1D4PHI1Z2n2_ME_L5L6_L1D4PHI1Z2),
.number_in2(VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2_number),
.read_add2(VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI1Z2_ME_L5L6_L1D4PHI1Z2),
.matchout(ME_L5L6_L1D4PHI1Z2_CM_L5L6_L1D4PHI1Z2),
.valid_data(ME_L5L6_L1D4PHI1Z2_CM_L5L6_L1D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D4PHI2Z1(
.number_in1(VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1_number),
.read_add1(VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1_read_add),
.vmstubin(VMS_L1D4PHI2Z1n4_ME_L5L6_L1D4PHI2Z1),
.number_in2(VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1_number),
.read_add2(VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI2Z1_ME_L5L6_L1D4PHI2Z1),
.matchout(ME_L5L6_L1D4PHI2Z1_CM_L5L6_L1D4PHI2Z1),
.valid_data(ME_L5L6_L1D4PHI2Z1_CM_L5L6_L1D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D4PHI2Z2(
.number_in1(VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2_number),
.read_add1(VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2_read_add),
.vmstubin(VMS_L1D4PHI2Z2n2_ME_L5L6_L1D4PHI2Z2),
.number_in2(VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2_number),
.read_add2(VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI2Z2_ME_L5L6_L1D4PHI2Z2),
.matchout(ME_L5L6_L1D4PHI2Z2_CM_L5L6_L1D4PHI2Z2),
.valid_data(ME_L5L6_L1D4PHI2Z2_CM_L5L6_L1D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D4PHI3Z1(
.number_in1(VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1_number),
.read_add1(VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1_read_add),
.vmstubin(VMS_L1D4PHI3Z1n4_ME_L5L6_L1D4PHI3Z1),
.number_in2(VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1_number),
.read_add2(VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI3Z1_ME_L5L6_L1D4PHI3Z1),
.matchout(ME_L5L6_L1D4PHI3Z1_CM_L5L6_L1D4PHI3Z1),
.valid_data(ME_L5L6_L1D4PHI3Z1_CM_L5L6_L1D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L1D4PHI3Z2(
.number_in1(VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2_number),
.read_add1(VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2_read_add),
.vmstubin(VMS_L1D4PHI3Z2n2_ME_L5L6_L1D4PHI3Z2),
.number_in2(VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2_number),
.read_add2(VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI3Z2_ME_L5L6_L1D4PHI3Z2),
.matchout(ME_L5L6_L1D4PHI3Z2_CM_L5L6_L1D4PHI3Z2),
.valid_data(ME_L5L6_L1D4PHI3Z2_CM_L5L6_L1D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D3PHI1Z1(
.number_in1(VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1_number),
.read_add1(VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1_read_add),
.vmstubin(VMS_L2D3PHI1Z1n3_ME_L5L6_L2D3PHI1Z1),
.number_in2(VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1_number),
.read_add2(VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI1Z1_ME_L5L6_L2D3PHI1Z1),
.matchout(ME_L5L6_L2D3PHI1Z1_CM_L5L6_L2D3PHI1Z1),
.valid_data(ME_L5L6_L2D3PHI1Z1_CM_L5L6_L2D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D3PHI1Z2(
.number_in1(VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2_number),
.read_add1(VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2_read_add),
.vmstubin(VMS_L2D3PHI1Z2n4_ME_L5L6_L2D3PHI1Z2),
.number_in2(VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2_number),
.read_add2(VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI1Z2_ME_L5L6_L2D3PHI1Z2),
.matchout(ME_L5L6_L2D3PHI1Z2_CM_L5L6_L2D3PHI1Z2),
.valid_data(ME_L5L6_L2D3PHI1Z2_CM_L5L6_L2D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D3PHI2Z1(
.number_in1(VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1_number),
.read_add1(VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1_read_add),
.vmstubin(VMS_L2D3PHI2Z1n4_ME_L5L6_L2D3PHI2Z1),
.number_in2(VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1_number),
.read_add2(VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI2Z1_ME_L5L6_L2D3PHI2Z1),
.matchout(ME_L5L6_L2D3PHI2Z1_CM_L5L6_L2D3PHI2Z1),
.valid_data(ME_L5L6_L2D3PHI2Z1_CM_L5L6_L2D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D3PHI2Z2(
.number_in1(VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2_number),
.read_add1(VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2_read_add),
.vmstubin(VMS_L2D3PHI2Z2n6_ME_L5L6_L2D3PHI2Z2),
.number_in2(VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2_number),
.read_add2(VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI2Z2_ME_L5L6_L2D3PHI2Z2),
.matchout(ME_L5L6_L2D3PHI2Z2_CM_L5L6_L2D3PHI2Z2),
.valid_data(ME_L5L6_L2D3PHI2Z2_CM_L5L6_L2D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D3PHI3Z1(
.number_in1(VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1_number),
.read_add1(VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1_read_add),
.vmstubin(VMS_L2D3PHI3Z1n4_ME_L5L6_L2D3PHI3Z1),
.number_in2(VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1_number),
.read_add2(VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI3Z1_ME_L5L6_L2D3PHI3Z1),
.matchout(ME_L5L6_L2D3PHI3Z1_CM_L5L6_L2D3PHI3Z1),
.valid_data(ME_L5L6_L2D3PHI3Z1_CM_L5L6_L2D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D3PHI3Z2(
.number_in1(VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2_number),
.read_add1(VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2_read_add),
.vmstubin(VMS_L2D3PHI3Z2n6_ME_L5L6_L2D3PHI3Z2),
.number_in2(VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2_number),
.read_add2(VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI3Z2_ME_L5L6_L2D3PHI3Z2),
.matchout(ME_L5L6_L2D3PHI3Z2_CM_L5L6_L2D3PHI3Z2),
.valid_data(ME_L5L6_L2D3PHI3Z2_CM_L5L6_L2D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D3PHI4Z1(
.number_in1(VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1_number),
.read_add1(VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1_read_add),
.vmstubin(VMS_L2D3PHI4Z1n3_ME_L5L6_L2D3PHI4Z1),
.number_in2(VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1_number),
.read_add2(VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI4Z1_ME_L5L6_L2D3PHI4Z1),
.matchout(ME_L5L6_L2D3PHI4Z1_CM_L5L6_L2D3PHI4Z1),
.valid_data(ME_L5L6_L2D3PHI4Z1_CM_L5L6_L2D3PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D3PHI4Z2(
.number_in1(VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2_number),
.read_add1(VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2_read_add),
.vmstubin(VMS_L2D3PHI4Z2n4_ME_L5L6_L2D3PHI4Z2),
.number_in2(VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2_number),
.read_add2(VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI4Z2_ME_L5L6_L2D3PHI4Z2),
.matchout(ME_L5L6_L2D3PHI4Z2_CM_L5L6_L2D3PHI4Z2),
.valid_data(ME_L5L6_L2D3PHI4Z2_CM_L5L6_L2D3PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D4PHI1Z1(
.number_in1(VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1_number),
.read_add1(VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1_read_add),
.vmstubin(VMS_L2D4PHI1Z1n4_ME_L5L6_L2D4PHI1Z1),
.number_in2(VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1_number),
.read_add2(VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI1Z1_ME_L5L6_L2D4PHI1Z1),
.matchout(ME_L5L6_L2D4PHI1Z1_CM_L5L6_L2D4PHI1Z1),
.valid_data(ME_L5L6_L2D4PHI1Z1_CM_L5L6_L2D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D4PHI1Z2(
.number_in1(VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2_number),
.read_add1(VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2_read_add),
.vmstubin(VMS_L2D4PHI1Z2n4_ME_L5L6_L2D4PHI1Z2),
.number_in2(VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2_number),
.read_add2(VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI1Z2_ME_L5L6_L2D4PHI1Z2),
.matchout(ME_L5L6_L2D4PHI1Z2_CM_L5L6_L2D4PHI1Z2),
.valid_data(ME_L5L6_L2D4PHI1Z2_CM_L5L6_L2D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D4PHI2Z1(
.number_in1(VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1_number),
.read_add1(VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1_read_add),
.vmstubin(VMS_L2D4PHI2Z1n6_ME_L5L6_L2D4PHI2Z1),
.number_in2(VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1_number),
.read_add2(VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI2Z1_ME_L5L6_L2D4PHI2Z1),
.matchout(ME_L5L6_L2D4PHI2Z1_CM_L5L6_L2D4PHI2Z1),
.valid_data(ME_L5L6_L2D4PHI2Z1_CM_L5L6_L2D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D4PHI2Z2(
.number_in1(VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2_number),
.read_add1(VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2_read_add),
.vmstubin(VMS_L2D4PHI2Z2n6_ME_L5L6_L2D4PHI2Z2),
.number_in2(VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2_number),
.read_add2(VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI2Z2_ME_L5L6_L2D4PHI2Z2),
.matchout(ME_L5L6_L2D4PHI2Z2_CM_L5L6_L2D4PHI2Z2),
.valid_data(ME_L5L6_L2D4PHI2Z2_CM_L5L6_L2D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D4PHI3Z1(
.number_in1(VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1_number),
.read_add1(VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1_read_add),
.vmstubin(VMS_L2D4PHI3Z1n6_ME_L5L6_L2D4PHI3Z1),
.number_in2(VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1_number),
.read_add2(VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI3Z1_ME_L5L6_L2D4PHI3Z1),
.matchout(ME_L5L6_L2D4PHI3Z1_CM_L5L6_L2D4PHI3Z1),
.valid_data(ME_L5L6_L2D4PHI3Z1_CM_L5L6_L2D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D4PHI3Z2(
.number_in1(VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2_number),
.read_add1(VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2_read_add),
.vmstubin(VMS_L2D4PHI3Z2n6_ME_L5L6_L2D4PHI3Z2),
.number_in2(VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2_number),
.read_add2(VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI3Z2_ME_L5L6_L2D4PHI3Z2),
.matchout(ME_L5L6_L2D4PHI3Z2_CM_L5L6_L2D4PHI3Z2),
.valid_data(ME_L5L6_L2D4PHI3Z2_CM_L5L6_L2D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D4PHI4Z1(
.number_in1(VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1_number),
.read_add1(VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1_read_add),
.vmstubin(VMS_L2D4PHI4Z1n4_ME_L5L6_L2D4PHI4Z1),
.number_in2(VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1_number),
.read_add2(VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI4Z1_ME_L5L6_L2D4PHI4Z1),
.matchout(ME_L5L6_L2D4PHI4Z1_CM_L5L6_L2D4PHI4Z1),
.valid_data(ME_L5L6_L2D4PHI4Z1_CM_L5L6_L2D4PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L2D4PHI4Z2(
.number_in1(VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2_number),
.read_add1(VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2_read_add),
.vmstubin(VMS_L2D4PHI4Z2n4_ME_L5L6_L2D4PHI4Z2),
.number_in2(VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2_number),
.read_add2(VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI4Z2_ME_L5L6_L2D4PHI4Z2),
.matchout(ME_L5L6_L2D4PHI4Z2_CM_L5L6_L2D4PHI4Z2),
.valid_data(ME_L5L6_L2D4PHI4Z2_CM_L5L6_L2D4PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D3PHI1Z1(
.number_in1(VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1_number),
.read_add1(VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1_read_add),
.vmstubin(VMS_L3D3PHI1Z1n6_ME_L5L6_L3D3PHI1Z1),
.number_in2(VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1_number),
.read_add2(VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI1Z1_ME_L5L6_L3D3PHI1Z1),
.matchout(ME_L5L6_L3D3PHI1Z1_CM_L5L6_L3D3PHI1Z1),
.valid_data(ME_L5L6_L3D3PHI1Z1_CM_L5L6_L3D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D3PHI1Z2(
.number_in1(VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2_number),
.read_add1(VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2_read_add),
.vmstubin(VMS_L3D3PHI1Z2n6_ME_L5L6_L3D3PHI1Z2),
.number_in2(VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2_number),
.read_add2(VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI1Z2_ME_L5L6_L3D3PHI1Z2),
.matchout(ME_L5L6_L3D3PHI1Z2_CM_L5L6_L3D3PHI1Z2),
.valid_data(ME_L5L6_L3D3PHI1Z2_CM_L5L6_L3D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D3PHI2Z1(
.number_in1(VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1_number),
.read_add1(VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1_read_add),
.vmstubin(VMS_L3D3PHI2Z1n6_ME_L5L6_L3D3PHI2Z1),
.number_in2(VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1_number),
.read_add2(VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI2Z1_ME_L5L6_L3D3PHI2Z1),
.matchout(ME_L5L6_L3D3PHI2Z1_CM_L5L6_L3D3PHI2Z1),
.valid_data(ME_L5L6_L3D3PHI2Z1_CM_L5L6_L3D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D3PHI2Z2(
.number_in1(VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2_number),
.read_add1(VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2_read_add),
.vmstubin(VMS_L3D3PHI2Z2n6_ME_L5L6_L3D3PHI2Z2),
.number_in2(VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2_number),
.read_add2(VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI2Z2_ME_L5L6_L3D3PHI2Z2),
.matchout(ME_L5L6_L3D3PHI2Z2_CM_L5L6_L3D3PHI2Z2),
.valid_data(ME_L5L6_L3D3PHI2Z2_CM_L5L6_L3D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D3PHI3Z1(
.number_in1(VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1_number),
.read_add1(VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1_read_add),
.vmstubin(VMS_L3D3PHI3Z1n6_ME_L5L6_L3D3PHI3Z1),
.number_in2(VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1_number),
.read_add2(VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI3Z1_ME_L5L6_L3D3PHI3Z1),
.matchout(ME_L5L6_L3D3PHI3Z1_CM_L5L6_L3D3PHI3Z1),
.valid_data(ME_L5L6_L3D3PHI3Z1_CM_L5L6_L3D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D3PHI3Z2(
.number_in1(VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2_number),
.read_add1(VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2_read_add),
.vmstubin(VMS_L3D3PHI3Z2n6_ME_L5L6_L3D3PHI3Z2),
.number_in2(VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2_number),
.read_add2(VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI3Z2_ME_L5L6_L3D3PHI3Z2),
.matchout(ME_L5L6_L3D3PHI3Z2_CM_L5L6_L3D3PHI3Z2),
.valid_data(ME_L5L6_L3D3PHI3Z2_CM_L5L6_L3D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D4PHI1Z1(
.number_in1(VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1_number),
.read_add1(VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1_read_add),
.vmstubin(VMS_L3D4PHI1Z1n6_ME_L5L6_L3D4PHI1Z1),
.number_in2(VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1_number),
.read_add2(VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI1Z1_ME_L5L6_L3D4PHI1Z1),
.matchout(ME_L5L6_L3D4PHI1Z1_CM_L5L6_L3D4PHI1Z1),
.valid_data(ME_L5L6_L3D4PHI1Z1_CM_L5L6_L3D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D4PHI1Z2(
.number_in1(VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2_number),
.read_add1(VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2_read_add),
.vmstubin(VMS_L3D4PHI1Z2n4_ME_L5L6_L3D4PHI1Z2),
.number_in2(VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2_number),
.read_add2(VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI1Z2_ME_L5L6_L3D4PHI1Z2),
.matchout(ME_L5L6_L3D4PHI1Z2_CM_L5L6_L3D4PHI1Z2),
.valid_data(ME_L5L6_L3D4PHI1Z2_CM_L5L6_L3D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D4PHI2Z1(
.number_in1(VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1_number),
.read_add1(VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1_read_add),
.vmstubin(VMS_L3D4PHI2Z1n6_ME_L5L6_L3D4PHI2Z1),
.number_in2(VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1_number),
.read_add2(VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI2Z1_ME_L5L6_L3D4PHI2Z1),
.matchout(ME_L5L6_L3D4PHI2Z1_CM_L5L6_L3D4PHI2Z1),
.valid_data(ME_L5L6_L3D4PHI2Z1_CM_L5L6_L3D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D4PHI2Z2(
.number_in1(VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2_number),
.read_add1(VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2_read_add),
.vmstubin(VMS_L3D4PHI2Z2n4_ME_L5L6_L3D4PHI2Z2),
.number_in2(VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2_number),
.read_add2(VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI2Z2_ME_L5L6_L3D4PHI2Z2),
.matchout(ME_L5L6_L3D4PHI2Z2_CM_L5L6_L3D4PHI2Z2),
.valid_data(ME_L5L6_L3D4PHI2Z2_CM_L5L6_L3D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D4PHI3Z1(
.number_in1(VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1_number),
.read_add1(VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1_read_add),
.vmstubin(VMS_L3D4PHI3Z1n6_ME_L5L6_L3D4PHI3Z1),
.number_in2(VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1_number),
.read_add2(VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI3Z1_ME_L5L6_L3D4PHI3Z1),
.matchout(ME_L5L6_L3D4PHI3Z1_CM_L5L6_L3D4PHI3Z1),
.valid_data(ME_L5L6_L3D4PHI3Z1_CM_L5L6_L3D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L3D4PHI3Z2(
.number_in1(VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2_number),
.read_add1(VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2_read_add),
.vmstubin(VMS_L3D4PHI3Z2n4_ME_L5L6_L3D4PHI3Z2),
.number_in2(VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2_number),
.read_add2(VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI3Z2_ME_L5L6_L3D4PHI3Z2),
.matchout(ME_L5L6_L3D4PHI3Z2_CM_L5L6_L3D4PHI3Z2),
.valid_data(ME_L5L6_L3D4PHI3Z2_CM_L5L6_L3D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D3PHI1Z1(
.number_in1(VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1_number),
.read_add1(VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1_read_add),
.vmstubin(VMS_L4D3PHI1Z1n3_ME_L5L6_L4D3PHI1Z1),
.number_in2(VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1_number),
.read_add2(VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI1Z1_ME_L5L6_L4D3PHI1Z1),
.matchout(ME_L5L6_L4D3PHI1Z1_CM_L5L6_L4D3PHI1Z1),
.valid_data(ME_L5L6_L4D3PHI1Z1_CM_L5L6_L4D3PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D3PHI1Z2(
.number_in1(VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2_number),
.read_add1(VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2_read_add),
.vmstubin(VMS_L4D3PHI1Z2n4_ME_L5L6_L4D3PHI1Z2),
.number_in2(VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2_number),
.read_add2(VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI1Z2_ME_L5L6_L4D3PHI1Z2),
.matchout(ME_L5L6_L4D3PHI1Z2_CM_L5L6_L4D3PHI1Z2),
.valid_data(ME_L5L6_L4D3PHI1Z2_CM_L5L6_L4D3PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D3PHI2Z1(
.number_in1(VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1_number),
.read_add1(VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1_read_add),
.vmstubin(VMS_L4D3PHI2Z1n4_ME_L5L6_L4D3PHI2Z1),
.number_in2(VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1_number),
.read_add2(VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI2Z1_ME_L5L6_L4D3PHI2Z1),
.matchout(ME_L5L6_L4D3PHI2Z1_CM_L5L6_L4D3PHI2Z1),
.valid_data(ME_L5L6_L4D3PHI2Z1_CM_L5L6_L4D3PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D3PHI2Z2(
.number_in1(VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2_number),
.read_add1(VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2_read_add),
.vmstubin(VMS_L4D3PHI2Z2n6_ME_L5L6_L4D3PHI2Z2),
.number_in2(VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2_number),
.read_add2(VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI2Z2_ME_L5L6_L4D3PHI2Z2),
.matchout(ME_L5L6_L4D3PHI2Z2_CM_L5L6_L4D3PHI2Z2),
.valid_data(ME_L5L6_L4D3PHI2Z2_CM_L5L6_L4D3PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D3PHI3Z1(
.number_in1(VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1_number),
.read_add1(VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1_read_add),
.vmstubin(VMS_L4D3PHI3Z1n4_ME_L5L6_L4D3PHI3Z1),
.number_in2(VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1_number),
.read_add2(VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI3Z1_ME_L5L6_L4D3PHI3Z1),
.matchout(ME_L5L6_L4D3PHI3Z1_CM_L5L6_L4D3PHI3Z1),
.valid_data(ME_L5L6_L4D3PHI3Z1_CM_L5L6_L4D3PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D3PHI3Z2(
.number_in1(VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2_number),
.read_add1(VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2_read_add),
.vmstubin(VMS_L4D3PHI3Z2n6_ME_L5L6_L4D3PHI3Z2),
.number_in2(VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2_number),
.read_add2(VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI3Z2_ME_L5L6_L4D3PHI3Z2),
.matchout(ME_L5L6_L4D3PHI3Z2_CM_L5L6_L4D3PHI3Z2),
.valid_data(ME_L5L6_L4D3PHI3Z2_CM_L5L6_L4D3PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D3PHI4Z1(
.number_in1(VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1_number),
.read_add1(VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1_read_add),
.vmstubin(VMS_L4D3PHI4Z1n3_ME_L5L6_L4D3PHI4Z1),
.number_in2(VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1_number),
.read_add2(VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI4Z1_ME_L5L6_L4D3PHI4Z1),
.matchout(ME_L5L6_L4D3PHI4Z1_CM_L5L6_L4D3PHI4Z1),
.valid_data(ME_L5L6_L4D3PHI4Z1_CM_L5L6_L4D3PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D3PHI4Z2(
.number_in1(VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2_number),
.read_add1(VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2_read_add),
.vmstubin(VMS_L4D3PHI4Z2n4_ME_L5L6_L4D3PHI4Z2),
.number_in2(VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2_number),
.read_add2(VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI4Z2_ME_L5L6_L4D3PHI4Z2),
.matchout(ME_L5L6_L4D3PHI4Z2_CM_L5L6_L4D3PHI4Z2),
.valid_data(ME_L5L6_L4D3PHI4Z2_CM_L5L6_L4D3PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D4PHI1Z1(
.number_in1(VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1_number),
.read_add1(VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1_read_add),
.vmstubin(VMS_L4D4PHI1Z1n4_ME_L5L6_L4D4PHI1Z1),
.number_in2(VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1_number),
.read_add2(VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI1Z1_ME_L5L6_L4D4PHI1Z1),
.matchout(ME_L5L6_L4D4PHI1Z1_CM_L5L6_L4D4PHI1Z1),
.valid_data(ME_L5L6_L4D4PHI1Z1_CM_L5L6_L4D4PHI1Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D4PHI1Z2(
.number_in1(VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2_number),
.read_add1(VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2_read_add),
.vmstubin(VMS_L4D4PHI1Z2n4_ME_L5L6_L4D4PHI1Z2),
.number_in2(VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2_number),
.read_add2(VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI1Z2_ME_L5L6_L4D4PHI1Z2),
.matchout(ME_L5L6_L4D4PHI1Z2_CM_L5L6_L4D4PHI1Z2),
.valid_data(ME_L5L6_L4D4PHI1Z2_CM_L5L6_L4D4PHI1Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D4PHI2Z1(
.number_in1(VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1_number),
.read_add1(VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1_read_add),
.vmstubin(VMS_L4D4PHI2Z1n6_ME_L5L6_L4D4PHI2Z1),
.number_in2(VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1_number),
.read_add2(VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI2Z1_ME_L5L6_L4D4PHI2Z1),
.matchout(ME_L5L6_L4D4PHI2Z1_CM_L5L6_L4D4PHI2Z1),
.valid_data(ME_L5L6_L4D4PHI2Z1_CM_L5L6_L4D4PHI2Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D4PHI2Z2(
.number_in1(VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2_number),
.read_add1(VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2_read_add),
.vmstubin(VMS_L4D4PHI2Z2n6_ME_L5L6_L4D4PHI2Z2),
.number_in2(VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2_number),
.read_add2(VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI2Z2_ME_L5L6_L4D4PHI2Z2),
.matchout(ME_L5L6_L4D4PHI2Z2_CM_L5L6_L4D4PHI2Z2),
.valid_data(ME_L5L6_L4D4PHI2Z2_CM_L5L6_L4D4PHI2Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D4PHI3Z1(
.number_in1(VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1_number),
.read_add1(VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1_read_add),
.vmstubin(VMS_L4D4PHI3Z1n6_ME_L5L6_L4D4PHI3Z1),
.number_in2(VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1_number),
.read_add2(VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI3Z1_ME_L5L6_L4D4PHI3Z1),
.matchout(ME_L5L6_L4D4PHI3Z1_CM_L5L6_L4D4PHI3Z1),
.valid_data(ME_L5L6_L4D4PHI3Z1_CM_L5L6_L4D4PHI3Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D4PHI3Z2(
.number_in1(VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2_number),
.read_add1(VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2_read_add),
.vmstubin(VMS_L4D4PHI3Z2n6_ME_L5L6_L4D4PHI3Z2),
.number_in2(VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2_number),
.read_add2(VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI3Z2_ME_L5L6_L4D4PHI3Z2),
.matchout(ME_L5L6_L4D4PHI3Z2_CM_L5L6_L4D4PHI3Z2),
.valid_data(ME_L5L6_L4D4PHI3Z2_CM_L5L6_L4D4PHI3Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D4PHI4Z1(
.number_in1(VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1_number),
.read_add1(VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1_read_add),
.vmstubin(VMS_L4D4PHI4Z1n4_ME_L5L6_L4D4PHI4Z1),
.number_in2(VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1_number),
.read_add2(VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI4Z1_ME_L5L6_L4D4PHI4Z1),
.matchout(ME_L5L6_L4D4PHI4Z1_CM_L5L6_L4D4PHI4Z1),
.valid_data(ME_L5L6_L4D4PHI4Z1_CM_L5L6_L4D4PHI4Z1_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchEngine  ME_L5L6_L4D4PHI4Z2(
.number_in1(VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2_number),
.read_add1(VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2_read_add),
.vmstubin(VMS_L4D4PHI4Z2n4_ME_L5L6_L4D4PHI4Z2),
.number_in2(VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2_number),
.read_add2(VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI4Z2_ME_L5L6_L4D4PHI4Z2),
.matchout(ME_L5L6_L4D4PHI4Z2_CM_L5L6_L4D4PHI4Z2),
.valid_data(ME_L5L6_L4D4PHI4Z2_CM_L5L6_L4D4PHI4Z2_wr_en),
.start(start7_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L1,`Z_L1,`R_L1,`PHID_L1,`ZD_L1,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L3L4_L1,`MC_z_L3L4_L1,`MC_zfactor_INNER) MC_L3L4_L1D3(
.number_in1(CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3_number),
.read_add1(CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3_read_add),
.match1in(CM_L3L4_L1D3PHI1Z1_MC_L3L4_L1D3),
.number_in2(CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3_number),
.read_add2(CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3_read_add),
.match2in(CM_L3L4_L1D3PHI1Z2_MC_L3L4_L1D3),
.number_in3(CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3_number),
.read_add3(CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3_read_add),
.match3in(CM_L3L4_L1D3PHI2Z1_MC_L3L4_L1D3),
.number_in4(CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3_number),
.read_add4(CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3_read_add),
.match4in(CM_L3L4_L1D3PHI2Z2_MC_L3L4_L1D3),
.number_in5(CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3_number),
.read_add5(CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3_read_add),
.match5in(CM_L3L4_L1D3PHI3Z1_MC_L3L4_L1D3),
.number_in6(CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3_number),
.read_add6(CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3_read_add),
.match6in(CM_L3L4_L1D3PHI3Z2_MC_L3L4_L1D3),
.read_add_allproj(AP_L3L4_L1D3_MC_L3L4_L1D3_read_add),
.allprojin(AP_L3L4_L1D3_MC_L3L4_L1D3),
.read_add_allstub(AS_L1D3n3_MC_L3L4_L1D3_read_add),
.allstubin(AS_L1D3n3_MC_L3L4_L1D3),
.matchoutminus(MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus),
.matchoutplus(MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus),
.matchout1(MC_L3L4_L1D3_FM_L3L4_L1D3),
.valid_matchminus(MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus_wr_en),
.valid_match(MC_L3L4_L1D3_FM_L3L4_L1D3_wr_en),
.start(start8_5),
.done(done8_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L1,`Z_L1,`R_L1,`PHID_L1,`ZD_L1,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L3L4_L1,`MC_z_L3L4_L1,`MC_zfactor_INNER) MC_L3L4_L1D4(
.number_in1(CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4_number),
.read_add1(CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4_read_add),
.match1in(CM_L3L4_L1D4PHI1Z1_MC_L3L4_L1D4),
.number_in2(CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4_number),
.read_add2(CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4_read_add),
.match2in(CM_L3L4_L1D4PHI1Z2_MC_L3L4_L1D4),
.number_in3(CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4_number),
.read_add3(CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4_read_add),
.match3in(CM_L3L4_L1D4PHI2Z1_MC_L3L4_L1D4),
.number_in4(CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4_number),
.read_add4(CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4_read_add),
.match4in(CM_L3L4_L1D4PHI2Z2_MC_L3L4_L1D4),
.number_in5(CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4_number),
.read_add5(CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4_read_add),
.match5in(CM_L3L4_L1D4PHI3Z1_MC_L3L4_L1D4),
.number_in6(CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4_number),
.read_add6(CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4_read_add),
.match6in(CM_L3L4_L1D4PHI3Z2_MC_L3L4_L1D4),
.read_add_allproj(AP_L3L4_L1D4_MC_L3L4_L1D4_read_add),
.allprojin(AP_L3L4_L1D4_MC_L3L4_L1D4),
.read_add_allstub(AS_L1D4n2_MC_L3L4_L1D4_read_add),
.allstubin(AS_L1D4n2_MC_L3L4_L1D4),
.matchoutminus(MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus),
.matchoutplus(MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus),
.matchout1(MC_L3L4_L1D4_FM_L3L4_L1D4),
.valid_matchminus(MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus_wr_en),
.valid_match(MC_L3L4_L1D4_FM_L3L4_L1D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L2,`Z_L2,`R_L2,`PHID_L2,`ZD_L2,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L3L4_L2,`MC_z_L3L4_L2,`MC_zfactor_INNER) MC_L3L4_L2D3(
.number_in1(CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3_number),
.read_add1(CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3_read_add),
.match1in(CM_L3L4_L2D3PHI1Z1_MC_L3L4_L2D3),
.number_in2(CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3_number),
.read_add2(CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3_read_add),
.match2in(CM_L3L4_L2D3PHI1Z2_MC_L3L4_L2D3),
.number_in3(CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3_number),
.read_add3(CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3_read_add),
.match3in(CM_L3L4_L2D3PHI2Z1_MC_L3L4_L2D3),
.number_in4(CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3_number),
.read_add4(CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3_read_add),
.match4in(CM_L3L4_L2D3PHI2Z2_MC_L3L4_L2D3),
.number_in5(CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3_number),
.read_add5(CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3_read_add),
.match5in(CM_L3L4_L2D3PHI3Z1_MC_L3L4_L2D3),
.number_in6(CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3_number),
.read_add6(CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3_read_add),
.match6in(CM_L3L4_L2D3PHI3Z2_MC_L3L4_L2D3),
.number_in7(CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3_number),
.read_add7(CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3_read_add),
.match7in(CM_L3L4_L2D3PHI4Z1_MC_L3L4_L2D3),
.number_in8(CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3_number),
.read_add8(CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3_read_add),
.match8in(CM_L3L4_L2D3PHI4Z2_MC_L3L4_L2D3),
.read_add_allproj(AP_L3L4_L2D3_MC_L3L4_L2D3_read_add),
.allprojin(AP_L3L4_L2D3_MC_L3L4_L2D3),
.read_add_allstub(AS_L2D3n2_MC_L3L4_L2D3_read_add),
.allstubin(AS_L2D3n2_MC_L3L4_L2D3),
.matchoutminus(MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus),
.matchoutplus(MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus),
.matchout1(MC_L3L4_L2D3_FM_L3L4_L2D3),
.valid_matchminus(MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus_wr_en),
.valid_match(MC_L3L4_L2D3_FM_L3L4_L2D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L2,`Z_L2,`R_L2,`PHID_L2,`ZD_L2,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L3L4_L2,`MC_z_L3L4_L2,`MC_zfactor_INNER) MC_L3L4_L2D4(
.number_in1(CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4_number),
.read_add1(CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4_read_add),
.match1in(CM_L3L4_L2D4PHI1Z1_MC_L3L4_L2D4),
.number_in2(CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4_number),
.read_add2(CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4_read_add),
.match2in(CM_L3L4_L2D4PHI1Z2_MC_L3L4_L2D4),
.number_in3(CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4_number),
.read_add3(CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4_read_add),
.match3in(CM_L3L4_L2D4PHI2Z1_MC_L3L4_L2D4),
.number_in4(CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4_number),
.read_add4(CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4_read_add),
.match4in(CM_L3L4_L2D4PHI2Z2_MC_L3L4_L2D4),
.number_in5(CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4_number),
.read_add5(CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4_read_add),
.match5in(CM_L3L4_L2D4PHI3Z1_MC_L3L4_L2D4),
.number_in6(CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4_number),
.read_add6(CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4_read_add),
.match6in(CM_L3L4_L2D4PHI3Z2_MC_L3L4_L2D4),
.number_in7(CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4_number),
.read_add7(CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4_read_add),
.match7in(CM_L3L4_L2D4PHI4Z1_MC_L3L4_L2D4),
.number_in8(CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4_number),
.read_add8(CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4_read_add),
.match8in(CM_L3L4_L2D4PHI4Z2_MC_L3L4_L2D4),
.read_add_allproj(AP_L3L4_L2D4_MC_L3L4_L2D4_read_add),
.allprojin(AP_L3L4_L2D4_MC_L3L4_L2D4),
.read_add_allstub(AS_L2D4n3_MC_L3L4_L2D4_read_add),
.allstubin(AS_L2D4n3_MC_L3L4_L2D4),
.matchoutminus(MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus),
.matchoutplus(MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus),
.matchout1(MC_L3L4_L2D4_FM_L3L4_L2D4),
.valid_matchminus(MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus_wr_en),
.valid_match(MC_L3L4_L2D4_FM_L3L4_L2D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L5,`Z_L5,`R_L5,`PHID_L5,`ZD_L5,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L3L4_L5,`MC_z_L3L4_L5,`MC_zfactor_OUTER) MC_L3L4_L5D3(
.number_in1(CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3_number),
.read_add1(CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3_read_add),
.match1in(CM_L3L4_L5D3PHI1Z1_MC_L3L4_L5D3),
.number_in2(CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3_number),
.read_add2(CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3_read_add),
.match2in(CM_L3L4_L5D3PHI1Z2_MC_L3L4_L5D3),
.number_in3(CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3_number),
.read_add3(CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3_read_add),
.match3in(CM_L3L4_L5D3PHI2Z1_MC_L3L4_L5D3),
.number_in4(CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3_number),
.read_add4(CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3_read_add),
.match4in(CM_L3L4_L5D3PHI2Z2_MC_L3L4_L5D3),
.number_in5(CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3_number),
.read_add5(CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3_read_add),
.match5in(CM_L3L4_L5D3PHI3Z1_MC_L3L4_L5D3),
.number_in6(CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3_number),
.read_add6(CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3_read_add),
.match6in(CM_L3L4_L5D3PHI3Z2_MC_L3L4_L5D3),
.read_add_allproj(AP_L3L4_L5D3_MC_L3L4_L5D3_read_add),
.allprojin(AP_L3L4_L5D3_MC_L3L4_L5D3),
.read_add_allstub(AS_L5D3n3_MC_L3L4_L5D3_read_add),
.allstubin(AS_L5D3n3_MC_L3L4_L5D3),
.matchoutminus(MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus),
.matchoutplus(MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus),
.matchout1(MC_L3L4_L5D3_FM_L3L4_L5D3),
.valid_matchminus(MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus_wr_en),
.valid_match(MC_L3L4_L5D3_FM_L3L4_L5D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L5,`Z_L5,`R_L5,`PHID_L5,`ZD_L5,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L3L4_L5,`MC_z_L3L4_L5,`MC_zfactor_OUTER) MC_L3L4_L5D4(
.number_in1(CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4_number),
.read_add1(CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4_read_add),
.match1in(CM_L3L4_L5D4PHI1Z1_MC_L3L4_L5D4),
.number_in2(CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4_number),
.read_add2(CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4_read_add),
.match2in(CM_L3L4_L5D4PHI1Z2_MC_L3L4_L5D4),
.number_in3(CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4_number),
.read_add3(CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4_read_add),
.match3in(CM_L3L4_L5D4PHI2Z1_MC_L3L4_L5D4),
.number_in4(CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4_number),
.read_add4(CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4_read_add),
.match4in(CM_L3L4_L5D4PHI2Z2_MC_L3L4_L5D4),
.number_in5(CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4_number),
.read_add5(CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4_read_add),
.match5in(CM_L3L4_L5D4PHI3Z1_MC_L3L4_L5D4),
.number_in6(CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4_number),
.read_add6(CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4_read_add),
.match6in(CM_L3L4_L5D4PHI3Z2_MC_L3L4_L5D4),
.read_add_allproj(AP_L3L4_L5D4_MC_L3L4_L5D4_read_add),
.allprojin(AP_L3L4_L5D4_MC_L3L4_L5D4),
.read_add_allstub(AS_L5D4n2_MC_L3L4_L5D4_read_add),
.allstubin(AS_L5D4n2_MC_L3L4_L5D4),
.matchoutminus(MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus),
.matchoutplus(MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus),
.matchout1(MC_L3L4_L5D4_FM_L3L4_L5D4),
.valid_matchminus(MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus_wr_en),
.valid_match(MC_L3L4_L5D4_FM_L3L4_L5D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L6,`Z_L6,`R_L6,`PHID_L6,`ZD_L6,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L3L4_L6,`MC_z_L3L4_L6,`MC_zfactor_OUTER) MC_L3L4_L6D3(
.number_in1(CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3_number),
.read_add1(CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3_read_add),
.match1in(CM_L3L4_L6D3PHI1Z1_MC_L3L4_L6D3),
.number_in2(CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3_number),
.read_add2(CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3_read_add),
.match2in(CM_L3L4_L6D3PHI1Z2_MC_L3L4_L6D3),
.number_in3(CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3_number),
.read_add3(CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3_read_add),
.match3in(CM_L3L4_L6D3PHI2Z1_MC_L3L4_L6D3),
.number_in4(CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3_number),
.read_add4(CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3_read_add),
.match4in(CM_L3L4_L6D3PHI2Z2_MC_L3L4_L6D3),
.number_in5(CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3_number),
.read_add5(CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3_read_add),
.match5in(CM_L3L4_L6D3PHI3Z1_MC_L3L4_L6D3),
.number_in6(CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3_number),
.read_add6(CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3_read_add),
.match6in(CM_L3L4_L6D3PHI3Z2_MC_L3L4_L6D3),
.number_in7(CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3_number),
.read_add7(CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3_read_add),
.match7in(CM_L3L4_L6D3PHI4Z1_MC_L3L4_L6D3),
.number_in8(CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3_number),
.read_add8(CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3_read_add),
.match8in(CM_L3L4_L6D3PHI4Z2_MC_L3L4_L6D3),
.read_add_allproj(AP_L3L4_L6D3_MC_L3L4_L6D3_read_add),
.allprojin(AP_L3L4_L6D3_MC_L3L4_L6D3),
.read_add_allstub(AS_L6D3n2_MC_L3L4_L6D3_read_add),
.allstubin(AS_L6D3n2_MC_L3L4_L6D3),
.matchoutminus(MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus),
.matchoutplus(MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus),
.matchout1(MC_L3L4_L6D3_FM_L3L4_L6D3),
.valid_matchminus(MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus_wr_en),
.valid_match(MC_L3L4_L6D3_FM_L3L4_L6D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L6,`Z_L6,`R_L6,`PHID_L6,`ZD_L6,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L3L4_L6,`MC_z_L3L4_L6,`MC_zfactor_OUTER) MC_L3L4_L6D4(
.number_in1(CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4_number),
.read_add1(CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4_read_add),
.match1in(CM_L3L4_L6D4PHI1Z1_MC_L3L4_L6D4),
.number_in2(CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4_number),
.read_add2(CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4_read_add),
.match2in(CM_L3L4_L6D4PHI1Z2_MC_L3L4_L6D4),
.number_in3(CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4_number),
.read_add3(CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4_read_add),
.match3in(CM_L3L4_L6D4PHI2Z1_MC_L3L4_L6D4),
.number_in4(CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4_number),
.read_add4(CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4_read_add),
.match4in(CM_L3L4_L6D4PHI2Z2_MC_L3L4_L6D4),
.number_in5(CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4_number),
.read_add5(CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4_read_add),
.match5in(CM_L3L4_L6D4PHI3Z1_MC_L3L4_L6D4),
.number_in6(CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4_number),
.read_add6(CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4_read_add),
.match6in(CM_L3L4_L6D4PHI3Z2_MC_L3L4_L6D4),
.number_in7(CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4_number),
.read_add7(CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4_read_add),
.match7in(CM_L3L4_L6D4PHI4Z1_MC_L3L4_L6D4),
.number_in8(CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4_number),
.read_add8(CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4_read_add),
.match8in(CM_L3L4_L6D4PHI4Z2_MC_L3L4_L6D4),
.read_add_allproj(AP_L3L4_L6D4_MC_L3L4_L6D4_read_add),
.allprojin(AP_L3L4_L6D4_MC_L3L4_L6D4),
.read_add_allstub(AS_L6D4n3_MC_L3L4_L6D4_read_add),
.allstubin(AS_L6D4n3_MC_L3L4_L6D4),
.matchoutminus(MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus),
.matchoutplus(MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus),
.matchout1(MC_L3L4_L6D4_FM_L3L4_L6D4),
.valid_matchminus(MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus_wr_en),
.valid_match(MC_L3L4_L6D4_FM_L3L4_L6D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator#(1'b1,`PHI_L1,`Z_L1,`R_L1,`PHID_L1,`ZD_L1,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L1,`MC_z_L5L6_L1,`MC_zfactor_INNER) MC_L5L6_L1D3(
.number_in1(CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3_number),
.read_add1(CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3_read_add),
.match1in(CM_L5L6_L1D3PHI1Z1_MC_L5L6_L1D3),
.number_in2(CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3_number),
.read_add2(CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3_read_add),
.match2in(CM_L5L6_L1D3PHI1Z2_MC_L5L6_L1D3),
.number_in3(CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3_number),
.read_add3(CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3_read_add),
.match3in(CM_L5L6_L1D3PHI2Z1_MC_L5L6_L1D3),
.number_in4(CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3_number),
.read_add4(CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3_read_add),
.match4in(CM_L5L6_L1D3PHI2Z2_MC_L5L6_L1D3),
.number_in5(CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3_number),
.read_add5(CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3_read_add),
.match5in(CM_L5L6_L1D3PHI3Z1_MC_L5L6_L1D3),
.number_in6(CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3_number),
.read_add6(CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3_read_add),
.match6in(CM_L5L6_L1D3PHI3Z2_MC_L5L6_L1D3),
.read_add_allproj(AP_L5L6_L1D3_MC_L5L6_L1D3_read_add),
.allprojin(AP_L5L6_L1D3_MC_L5L6_L1D3),
.read_add_allstub(AS_L1D3n4_MC_L5L6_L1D3_read_add),
.allstubin(AS_L1D3n4_MC_L5L6_L1D3),
.matchoutminus(MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus),
.matchoutplus(MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus),
.matchout1(MC_L5L6_L1D3_FM_L5L6_L1D3),
.valid_matchminus(MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus_wr_en),
.valid_match(MC_L5L6_L1D3_FM_L5L6_L1D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L1,`Z_L1,`R_L1,`PHID_L1,`ZD_L1,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L1,`MC_z_L5L6_L1,`MC_zfactor_INNER) MC_L5L6_L1D4(
.number_in1(CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4_number),
.read_add1(CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4_read_add),
.match1in(CM_L5L6_L1D4PHI1Z1_MC_L5L6_L1D4),
.number_in2(CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4_number),
.read_add2(CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4_read_add),
.match2in(CM_L5L6_L1D4PHI1Z2_MC_L5L6_L1D4),
.number_in3(CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4_number),
.read_add3(CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4_read_add),
.match3in(CM_L5L6_L1D4PHI2Z1_MC_L5L6_L1D4),
.number_in4(CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4_number),
.read_add4(CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4_read_add),
.match4in(CM_L5L6_L1D4PHI2Z2_MC_L5L6_L1D4),
.number_in5(CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4_number),
.read_add5(CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4_read_add),
.match5in(CM_L5L6_L1D4PHI3Z1_MC_L5L6_L1D4),
.number_in6(CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4_number),
.read_add6(CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4_read_add),
.match6in(CM_L5L6_L1D4PHI3Z2_MC_L5L6_L1D4),
.read_add_allproj(AP_L5L6_L1D4_MC_L5L6_L1D4_read_add),
.allprojin(AP_L5L6_L1D4_MC_L5L6_L1D4),
.read_add_allstub(AS_L1D4n3_MC_L5L6_L1D4_read_add),
.allstubin(AS_L1D4n3_MC_L5L6_L1D4),
.matchoutminus(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus),
.matchoutplus(MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus),
.matchout1(MC_L5L6_L1D4_FM_L5L6_L1D4),
.valid_matchminus(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus_wr_en),
.valid_match(MC_L5L6_L1D4_FM_L5L6_L1D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L2,`Z_L2,`R_L2,`PHID_L2,`ZD_L2,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L2,`MC_z_L5L6_L2,`MC_zfactor_INNER) MC_L5L6_L2D3(
.number_in1(CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3_number),
.read_add1(CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3_read_add),
.match1in(CM_L5L6_L2D3PHI1Z1_MC_L5L6_L2D3),
.number_in2(CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3_number),
.read_add2(CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3_read_add),
.match2in(CM_L5L6_L2D3PHI1Z2_MC_L5L6_L2D3),
.number_in3(CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3_number),
.read_add3(CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3_read_add),
.match3in(CM_L5L6_L2D3PHI2Z1_MC_L5L6_L2D3),
.number_in4(CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3_number),
.read_add4(CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3_read_add),
.match4in(CM_L5L6_L2D3PHI2Z2_MC_L5L6_L2D3),
.number_in5(CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3_number),
.read_add5(CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3_read_add),
.match5in(CM_L5L6_L2D3PHI3Z1_MC_L5L6_L2D3),
.number_in6(CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3_number),
.read_add6(CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3_read_add),
.match6in(CM_L5L6_L2D3PHI3Z2_MC_L5L6_L2D3),
.number_in7(CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3_number),
.read_add7(CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3_read_add),
.match7in(CM_L5L6_L2D3PHI4Z1_MC_L5L6_L2D3),
.number_in8(CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3_number),
.read_add8(CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3_read_add),
.match8in(CM_L5L6_L2D3PHI4Z2_MC_L5L6_L2D3),
.read_add_allproj(AP_L5L6_L2D3_MC_L5L6_L2D3_read_add),
.allprojin(AP_L5L6_L2D3_MC_L5L6_L2D3),
.read_add_allstub(AS_L2D3n3_MC_L5L6_L2D3_read_add),
.allstubin(AS_L2D3n3_MC_L5L6_L2D3),
.matchoutminus(MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus),
.matchoutplus(MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus),
.matchout1(MC_L5L6_L2D3_FM_L5L6_L2D3),
.valid_matchminus(MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus_wr_en),
.valid_match(MC_L5L6_L2D3_FM_L5L6_L2D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L2,`Z_L2,`R_L2,`PHID_L2,`ZD_L2,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L2,`MC_z_L5L6_L2,`MC_zfactor_INNER) MC_L5L6_L2D4(
.number_in1(CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4_number),
.read_add1(CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4_read_add),
.match1in(CM_L5L6_L2D4PHI1Z1_MC_L5L6_L2D4),
.number_in2(CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4_number),
.read_add2(CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4_read_add),
.match2in(CM_L5L6_L2D4PHI1Z2_MC_L5L6_L2D4),
.number_in3(CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4_number),
.read_add3(CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4_read_add),
.match3in(CM_L5L6_L2D4PHI2Z1_MC_L5L6_L2D4),
.number_in4(CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4_number),
.read_add4(CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4_read_add),
.match4in(CM_L5L6_L2D4PHI2Z2_MC_L5L6_L2D4),
.number_in5(CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4_number),
.read_add5(CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4_read_add),
.match5in(CM_L5L6_L2D4PHI3Z1_MC_L5L6_L2D4),
.number_in6(CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4_number),
.read_add6(CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4_read_add),
.match6in(CM_L5L6_L2D4PHI3Z2_MC_L5L6_L2D4),
.number_in7(CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4_number),
.read_add7(CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4_read_add),
.match7in(CM_L5L6_L2D4PHI4Z1_MC_L5L6_L2D4),
.number_in8(CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4_number),
.read_add8(CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4_read_add),
.match8in(CM_L5L6_L2D4PHI4Z2_MC_L5L6_L2D4),
.read_add_allproj(AP_L5L6_L2D4_MC_L5L6_L2D4_read_add),
.allprojin(AP_L5L6_L2D4_MC_L5L6_L2D4),
.read_add_allstub(AS_L2D4n4_MC_L5L6_L2D4_read_add),
.allstubin(AS_L2D4n4_MC_L5L6_L2D4),
.matchoutminus(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus),
.matchoutplus(MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus),
.matchout1(MC_L5L6_L2D4_FM_L5L6_L2D4),
.valid_matchminus(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus_wr_en),
.valid_match(MC_L5L6_L2D4_FM_L5L6_L2D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L3,`Z_L3,`R_L3,`PHID_L3,`ZD_L3,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L3,`MC_z_L5L6_L3,`MC_zfactor_INNER) MC_L5L6_L3D3(
.number_in1(CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3_number),
.read_add1(CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3_read_add),
.match1in(CM_L5L6_L3D3PHI1Z1_MC_L5L6_L3D3),
.number_in2(CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3_number),
.read_add2(CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3_read_add),
.match2in(CM_L5L6_L3D3PHI1Z2_MC_L5L6_L3D3),
.number_in3(CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3_number),
.read_add3(CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3_read_add),
.match3in(CM_L5L6_L3D3PHI2Z1_MC_L5L6_L3D3),
.number_in4(CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3_number),
.read_add4(CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3_read_add),
.match4in(CM_L5L6_L3D3PHI2Z2_MC_L5L6_L3D3),
.number_in5(CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3_number),
.read_add5(CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3_read_add),
.match5in(CM_L5L6_L3D3PHI3Z1_MC_L5L6_L3D3),
.number_in6(CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3_number),
.read_add6(CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3_read_add),
.match6in(CM_L5L6_L3D3PHI3Z2_MC_L5L6_L3D3),
.read_add_allproj(AP_L5L6_L3D3_MC_L5L6_L3D3_read_add),
.allprojin(AP_L5L6_L3D3_MC_L5L6_L3D3),
.read_add_allstub(AS_L3D3n3_MC_L5L6_L3D3_read_add),
.allstubin(AS_L3D3n3_MC_L5L6_L3D3),
.matchoutminus(MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus),
.matchoutplus(MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus),
.matchout1(MC_L5L6_L3D3_FM_L5L6_L3D3),
.valid_matchminus(MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus_wr_en),
.valid_match(MC_L5L6_L3D3_FM_L5L6_L3D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L3,`Z_L3,`R_L3,`PHID_L3,`ZD_L3,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L3,`MC_z_L5L6_L3,`MC_zfactor_INNER) MC_L5L6_L3D4(
.number_in1(CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4_number),
.read_add1(CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4_read_add),
.match1in(CM_L5L6_L3D4PHI1Z1_MC_L5L6_L3D4),
.number_in2(CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4_number),
.read_add2(CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4_read_add),
.match2in(CM_L5L6_L3D4PHI1Z2_MC_L5L6_L3D4),
.number_in3(CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4_number),
.read_add3(CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4_read_add),
.match3in(CM_L5L6_L3D4PHI2Z1_MC_L5L6_L3D4),
.number_in4(CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4_number),
.read_add4(CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4_read_add),
.match4in(CM_L5L6_L3D4PHI2Z2_MC_L5L6_L3D4),
.number_in5(CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4_number),
.read_add5(CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4_read_add),
.match5in(CM_L5L6_L3D4PHI3Z1_MC_L5L6_L3D4),
.number_in6(CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4_number),
.read_add6(CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4_read_add),
.match6in(CM_L5L6_L3D4PHI3Z2_MC_L5L6_L3D4),
.read_add_allproj(AP_L5L6_L3D4_MC_L5L6_L3D4_read_add),
.allprojin(AP_L5L6_L3D4_MC_L5L6_L3D4),
.read_add_allstub(AS_L3D4n2_MC_L5L6_L3D4_read_add),
.allstubin(AS_L3D4n2_MC_L5L6_L3D4),
.matchoutminus(MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus),
.matchoutplus(MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus),
.matchout1(MC_L5L6_L3D4_FM_L5L6_L3D4),
.valid_matchminus(MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus_wr_en),
.valid_match(MC_L5L6_L3D4_FM_L5L6_L3D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L4,`Z_L4,`R_L4,`PHID_L4,`ZD_L4,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L5L6_L4,`MC_z_L5L6_L4,`MC_zfactor_OUTER) MC_L5L6_L4D3(
.number_in1(CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3_number),
.read_add1(CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3_read_add),
.match1in(CM_L5L6_L4D3PHI1Z1_MC_L5L6_L4D3),
.number_in2(CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3_number),
.read_add2(CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3_read_add),
.match2in(CM_L5L6_L4D3PHI1Z2_MC_L5L6_L4D3),
.number_in3(CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3_number),
.read_add3(CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3_read_add),
.match3in(CM_L5L6_L4D3PHI2Z1_MC_L5L6_L4D3),
.number_in4(CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3_number),
.read_add4(CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3_read_add),
.match4in(CM_L5L6_L4D3PHI2Z2_MC_L5L6_L4D3),
.number_in5(CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3_number),
.read_add5(CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3_read_add),
.match5in(CM_L5L6_L4D3PHI3Z1_MC_L5L6_L4D3),
.number_in6(CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3_number),
.read_add6(CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3_read_add),
.match6in(CM_L5L6_L4D3PHI3Z2_MC_L5L6_L4D3),
.number_in7(CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3_number),
.read_add7(CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3_read_add),
.match7in(CM_L5L6_L4D3PHI4Z1_MC_L5L6_L4D3),
.number_in8(CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3_number),
.read_add8(CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3_read_add),
.match8in(CM_L5L6_L4D3PHI4Z2_MC_L5L6_L4D3),
.read_add_allproj(AP_L5L6_L4D3_MC_L5L6_L4D3_read_add),
.allprojin(AP_L5L6_L4D3_MC_L5L6_L4D3),
.read_add_allstub(AS_L4D3n2_MC_L5L6_L4D3_read_add),
.allstubin(AS_L4D3n2_MC_L5L6_L4D3),
.matchoutminus(MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus),
.matchoutplus(MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus),
.matchout1(MC_L5L6_L4D3_FM_L5L6_L4D3),
.valid_matchminus(MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus_wr_en),
.valid_match(MC_L5L6_L4D3_FM_L5L6_L4D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L4,`Z_L4,`R_L4,`PHID_L4,`ZD_L4,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L5L6_L4,`MC_z_L5L6_L4,`MC_zfactor_OUTER) MC_L5L6_L4D4(
.number_in1(CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4_number),
.read_add1(CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4_read_add),
.match1in(CM_L5L6_L4D4PHI1Z1_MC_L5L6_L4D4),
.number_in2(CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4_number),
.read_add2(CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4_read_add),
.match2in(CM_L5L6_L4D4PHI1Z2_MC_L5L6_L4D4),
.number_in3(CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4_number),
.read_add3(CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4_read_add),
.match3in(CM_L5L6_L4D4PHI2Z1_MC_L5L6_L4D4),
.number_in4(CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4_number),
.read_add4(CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4_read_add),
.match4in(CM_L5L6_L4D4PHI2Z2_MC_L5L6_L4D4),
.number_in5(CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4_number),
.read_add5(CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4_read_add),
.match5in(CM_L5L6_L4D4PHI3Z1_MC_L5L6_L4D4),
.number_in6(CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4_number),
.read_add6(CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4_read_add),
.match6in(CM_L5L6_L4D4PHI3Z2_MC_L5L6_L4D4),
.number_in7(CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4_number),
.read_add7(CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4_read_add),
.match7in(CM_L5L6_L4D4PHI4Z1_MC_L5L6_L4D4),
.number_in8(CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4_number),
.read_add8(CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4_read_add),
.match8in(CM_L5L6_L4D4PHI4Z2_MC_L5L6_L4D4),
.read_add_allproj(AP_L5L6_L4D4_MC_L5L6_L4D4_read_add),
.allprojin(AP_L5L6_L4D4_MC_L5L6_L4D4),
.read_add_allstub(AS_L4D4n3_MC_L5L6_L4D4_read_add),
.allstubin(AS_L4D4n3_MC_L5L6_L4D4),
.matchoutminus(MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus),
.matchoutplus(MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus),
.matchout1(MC_L5L6_L4D4_FM_L5L6_L4D4),
.valid_matchminus(MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus_wr_en),
.valid_match(MC_L5L6_L4D4_FM_L5L6_L4D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L3,`Z_L3,`R_L3,`PHID_L3,`ZD_L3,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L1L2_L3,`MC_z_L1L2_L3,`MC_zfactor_INNER) MC_L1L2_L3D3(
.number_in1(CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3_number),
.read_add1(CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3_read_add),
.match1in(CM_L1L2_L3D3PHI1Z1_MC_L1L2_L3D3),
.number_in2(CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3_number),
.read_add2(CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3_read_add),
.match2in(CM_L1L2_L3D3PHI1Z2_MC_L1L2_L3D3),
.number_in3(CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3_number),
.read_add3(CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3_read_add),
.match3in(CM_L1L2_L3D3PHI2Z1_MC_L1L2_L3D3),
.number_in4(CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3_number),
.read_add4(CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3_read_add),
.match4in(CM_L1L2_L3D3PHI2Z2_MC_L1L2_L3D3),
.number_in5(CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3_number),
.read_add5(CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3_read_add),
.match5in(CM_L1L2_L3D3PHI3Z1_MC_L1L2_L3D3),
.number_in6(CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3_number),
.read_add6(CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3_read_add),
.match6in(CM_L1L2_L3D3PHI3Z2_MC_L1L2_L3D3),
.read_add_allproj(AP_L1L2_L3D3_MC_L1L2_L3D3_read_add),
.allprojin(AP_L1L2_L3D3_MC_L1L2_L3D3),
.read_add_allstub(AS_L3D3n4_MC_L1L2_L3D3_read_add),
.allstubin(AS_L3D3n4_MC_L1L2_L3D3),
.matchoutminus(MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus),
.matchoutplus(MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus),
.matchout1(MC_L1L2_L3D3_FM_L1L2_L3D3),
.valid_matchminus(MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus_wr_en),
.valid_match(MC_L1L2_L3D3_FM_L1L2_L3D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b1,`PHI_L3,`Z_L3,`R_L3,`PHID_L3,`ZD_L3,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L1L2_L3,`MC_z_L1L2_L3,`MC_zfactor_INNER) MC_L1L2_L3D4(
.number_in1(CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4_number),
.read_add1(CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4_read_add),
.match1in(CM_L1L2_L3D4PHI1Z1_MC_L1L2_L3D4),
.number_in2(CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4_number),
.read_add2(CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4_read_add),
.match2in(CM_L1L2_L3D4PHI1Z2_MC_L1L2_L3D4),
.number_in3(CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4_number),
.read_add3(CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4_read_add),
.match3in(CM_L1L2_L3D4PHI2Z1_MC_L1L2_L3D4),
.number_in4(CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4_number),
.read_add4(CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4_read_add),
.match4in(CM_L1L2_L3D4PHI2Z2_MC_L1L2_L3D4),
.number_in5(CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4_number),
.read_add5(CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4_read_add),
.match5in(CM_L1L2_L3D4PHI3Z1_MC_L1L2_L3D4),
.number_in6(CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4_number),
.read_add6(CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4_read_add),
.match6in(CM_L1L2_L3D4PHI3Z2_MC_L1L2_L3D4),
.read_add_allproj(AP_L1L2_L3D4_MC_L1L2_L3D4_read_add),
.allprojin(AP_L1L2_L3D4_MC_L1L2_L3D4),
.read_add_allstub(AS_L3D4n3_MC_L1L2_L3D4_read_add),
.allstubin(AS_L3D4n3_MC_L1L2_L3D4),
.matchoutminus(MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus),
.matchoutplus(MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus),
.matchout1(MC_L1L2_L3D4_FM_L1L2_L3D4),
.valid_matchminus(MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus_wr_en),
.valid_match(MC_L1L2_L3D4_FM_L1L2_L3D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L4,`Z_L4,`R_L4,`PHID_L4,`ZD_L4,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L4,`MC_z_L1L2_L4,`MC_zfactor_OUTER) MC_L1L2_L4D3(
.number_in1(CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3_number),
.read_add1(CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3_read_add),
.match1in(CM_L1L2_L4D3PHI1Z1_MC_L1L2_L4D3),
.number_in2(CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3_number),
.read_add2(CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3_read_add),
.match2in(CM_L1L2_L4D3PHI1Z2_MC_L1L2_L4D3),
.number_in3(CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3_number),
.read_add3(CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3_read_add),
.match3in(CM_L1L2_L4D3PHI2Z1_MC_L1L2_L4D3),
.number_in4(CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3_number),
.read_add4(CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3_read_add),
.match4in(CM_L1L2_L4D3PHI2Z2_MC_L1L2_L4D3),
.number_in5(CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3_number),
.read_add5(CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3_read_add),
.match5in(CM_L1L2_L4D3PHI3Z1_MC_L1L2_L4D3),
.number_in6(CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3_number),
.read_add6(CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3_read_add),
.match6in(CM_L1L2_L4D3PHI3Z2_MC_L1L2_L4D3),
.number_in7(CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3_number),
.read_add7(CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3_read_add),
.match7in(CM_L1L2_L4D3PHI4Z1_MC_L1L2_L4D3),
.number_in8(CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3_number),
.read_add8(CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3_read_add),
.match8in(CM_L1L2_L4D3PHI4Z2_MC_L1L2_L4D3),
.read_add_allproj(AP_L1L2_L4D3_MC_L1L2_L4D3_read_add),
.allprojin(AP_L1L2_L4D3_MC_L1L2_L4D3),
.read_add_allstub(AS_L4D3n3_MC_L1L2_L4D3_read_add),
.allstubin(AS_L4D3n3_MC_L1L2_L4D3),
.matchoutminus(MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus),
.matchoutplus(MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus),
.matchout1(MC_L1L2_L4D3_FM_L1L2_L4D3),
.valid_matchminus(MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus_wr_en),
.valid_match(MC_L1L2_L4D3_FM_L1L2_L4D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L4,`Z_L4,`R_L4,`PHID_L4,`ZD_L4,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L4,`MC_z_L1L2_L4,`MC_zfactor_OUTER) MC_L1L2_L4D4(
.number_in1(CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4_number),
.read_add1(CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4_read_add),
.match1in(CM_L1L2_L4D4PHI1Z1_MC_L1L2_L4D4),
.number_in2(CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4_number),
.read_add2(CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4_read_add),
.match2in(CM_L1L2_L4D4PHI1Z2_MC_L1L2_L4D4),
.number_in3(CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4_number),
.read_add3(CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4_read_add),
.match3in(CM_L1L2_L4D4PHI2Z1_MC_L1L2_L4D4),
.number_in4(CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4_number),
.read_add4(CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4_read_add),
.match4in(CM_L1L2_L4D4PHI2Z2_MC_L1L2_L4D4),
.number_in5(CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4_number),
.read_add5(CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4_read_add),
.match5in(CM_L1L2_L4D4PHI3Z1_MC_L1L2_L4D4),
.number_in6(CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4_number),
.read_add6(CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4_read_add),
.match6in(CM_L1L2_L4D4PHI3Z2_MC_L1L2_L4D4),
.number_in7(CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4_number),
.read_add7(CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4_read_add),
.match7in(CM_L1L2_L4D4PHI4Z1_MC_L1L2_L4D4),
.number_in8(CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4_number),
.read_add8(CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4_read_add),
.match8in(CM_L1L2_L4D4PHI4Z2_MC_L1L2_L4D4),
.read_add_allproj(AP_L1L2_L4D4_MC_L1L2_L4D4_read_add),
.allprojin(AP_L1L2_L4D4_MC_L1L2_L4D4),
.read_add_allstub(AS_L4D4n4_MC_L1L2_L4D4_read_add),
.allstubin(AS_L4D4n4_MC_L1L2_L4D4),
.matchoutminus(MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus),
.matchoutplus(MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus),
.matchout1(MC_L1L2_L4D4_FM_L1L2_L4D4),
.valid_matchminus(MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus_wr_en),
.valid_match(MC_L1L2_L4D4_FM_L1L2_L4D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L5,`Z_L5,`R_L5,`PHID_L5,`ZD_L5,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L5,`MC_z_L1L2_L5,`MC_zfactor_OUTER) MC_L1L2_L5D3(
.number_in1(CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3_number),
.read_add1(CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3_read_add),
.match1in(CM_L1L2_L5D3PHI1Z1_MC_L1L2_L5D3),
.number_in2(CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3_number),
.read_add2(CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3_read_add),
.match2in(CM_L1L2_L5D3PHI1Z2_MC_L1L2_L5D3),
.number_in3(CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3_number),
.read_add3(CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3_read_add),
.match3in(CM_L1L2_L5D3PHI2Z1_MC_L1L2_L5D3),
.number_in4(CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3_number),
.read_add4(CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3_read_add),
.match4in(CM_L1L2_L5D3PHI2Z2_MC_L1L2_L5D3),
.number_in5(CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3_number),
.read_add5(CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3_read_add),
.match5in(CM_L1L2_L5D3PHI3Z1_MC_L1L2_L5D3),
.number_in6(CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3_number),
.read_add6(CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3_read_add),
.match6in(CM_L1L2_L5D3PHI3Z2_MC_L1L2_L5D3),
.read_add_allproj(AP_L1L2_L5D3_MC_L1L2_L5D3_read_add),
.allprojin(AP_L1L2_L5D3_MC_L1L2_L5D3),
.read_add_allstub(AS_L5D3n4_MC_L1L2_L5D3_read_add),
.allstubin(AS_L5D3n4_MC_L1L2_L5D3),
.matchoutminus(MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus),
.matchoutplus(MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus),
.matchout1(MC_L1L2_L5D3_FM_L1L2_L5D3),
.valid_matchminus(MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus_wr_en),
.valid_match(MC_L1L2_L5D3_FM_L1L2_L5D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L5,`Z_L5,`R_L5,`PHID_L5,`ZD_L5,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L5,`MC_z_L1L2_L5,`MC_zfactor_OUTER) MC_L1L2_L5D4(
.number_in1(CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4_number),
.read_add1(CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4_read_add),
.match1in(CM_L1L2_L5D4PHI1Z1_MC_L1L2_L5D4),
.number_in2(CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4_number),
.read_add2(CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4_read_add),
.match2in(CM_L1L2_L5D4PHI1Z2_MC_L1L2_L5D4),
.number_in3(CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4_number),
.read_add3(CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4_read_add),
.match3in(CM_L1L2_L5D4PHI2Z1_MC_L1L2_L5D4),
.number_in4(CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4_number),
.read_add4(CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4_read_add),
.match4in(CM_L1L2_L5D4PHI2Z2_MC_L1L2_L5D4),
.number_in5(CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4_number),
.read_add5(CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4_read_add),
.match5in(CM_L1L2_L5D4PHI3Z1_MC_L1L2_L5D4),
.number_in6(CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4_number),
.read_add6(CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4_read_add),
.match6in(CM_L1L2_L5D4PHI3Z2_MC_L1L2_L5D4),
.read_add_allproj(AP_L1L2_L5D4_MC_L1L2_L5D4_read_add),
.allprojin(AP_L1L2_L5D4_MC_L1L2_L5D4),
.read_add_allstub(AS_L5D4n3_MC_L1L2_L5D4_read_add),
.allstubin(AS_L5D4n3_MC_L1L2_L5D4),
.matchoutminus(MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus),
.matchoutplus(MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus),
.matchout1(MC_L1L2_L5D4_FM_L1L2_L5D4),
.valid_matchminus(MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus_wr_en),
.valid_match(MC_L1L2_L5D4_FM_L1L2_L5D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L6,`Z_L6,`R_L6,`PHID_L6,`ZD_L6,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L6,`MC_z_L1L2_L6,`MC_zfactor_OUTER) MC_L1L2_L6D3(
.number_in1(CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3_number),
.read_add1(CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3_read_add),
.match1in(CM_L1L2_L6D3PHI1Z1_MC_L1L2_L6D3),
.number_in2(CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3_number),
.read_add2(CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3_read_add),
.match2in(CM_L1L2_L6D3PHI1Z2_MC_L1L2_L6D3),
.number_in3(CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3_number),
.read_add3(CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3_read_add),
.match3in(CM_L1L2_L6D3PHI2Z1_MC_L1L2_L6D3),
.number_in4(CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3_number),
.read_add4(CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3_read_add),
.match4in(CM_L1L2_L6D3PHI2Z2_MC_L1L2_L6D3),
.number_in5(CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3_number),
.read_add5(CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3_read_add),
.match5in(CM_L1L2_L6D3PHI3Z1_MC_L1L2_L6D3),
.number_in6(CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3_number),
.read_add6(CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3_read_add),
.match6in(CM_L1L2_L6D3PHI3Z2_MC_L1L2_L6D3),
.number_in7(CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3_number),
.read_add7(CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3_read_add),
.match7in(CM_L1L2_L6D3PHI4Z1_MC_L1L2_L6D3),
.number_in8(CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3_number),
.read_add8(CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3_read_add),
.match8in(CM_L1L2_L6D3PHI4Z2_MC_L1L2_L6D3),
.read_add_allproj(AP_L1L2_L6D3_MC_L1L2_L6D3_read_add),
.allprojin(AP_L1L2_L6D3_MC_L1L2_L6D3),
.read_add_allstub(AS_L6D3n3_MC_L1L2_L6D3_read_add),
.allstubin(AS_L6D3n3_MC_L1L2_L6D3),
.matchoutminus(MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus),
.matchoutplus(MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus),
.matchout1(MC_L1L2_L6D3_FM_L1L2_L6D3),
.valid_matchminus(MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus_wr_en),
.valid_match(MC_L1L2_L6D3_FM_L1L2_L6D3_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchCalculator #(1'b0,`PHI_L6,`Z_L6,`R_L6,`PHID_L6,`ZD_L6,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L6,`MC_z_L1L2_L6,`MC_zfactor_OUTER) MC_L1L2_L6D4(
.number_in1(CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4_number),
.read_add1(CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4_read_add),
.match1in(CM_L1L2_L6D4PHI1Z1_MC_L1L2_L6D4),
.number_in2(CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4_number),
.read_add2(CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4_read_add),
.match2in(CM_L1L2_L6D4PHI1Z2_MC_L1L2_L6D4),
.number_in3(CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4_number),
.read_add3(CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4_read_add),
.match3in(CM_L1L2_L6D4PHI2Z1_MC_L1L2_L6D4),
.number_in4(CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4_number),
.read_add4(CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4_read_add),
.match4in(CM_L1L2_L6D4PHI2Z2_MC_L1L2_L6D4),
.number_in5(CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4_number),
.read_add5(CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4_read_add),
.match5in(CM_L1L2_L6D4PHI3Z1_MC_L1L2_L6D4),
.number_in6(CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4_number),
.read_add6(CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4_read_add),
.match6in(CM_L1L2_L6D4PHI3Z2_MC_L1L2_L6D4),
.number_in7(CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4_number),
.read_add7(CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4_read_add),
.match7in(CM_L1L2_L6D4PHI4Z1_MC_L1L2_L6D4),
.number_in8(CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4_number),
.read_add8(CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4_read_add),
.match8in(CM_L1L2_L6D4PHI4Z2_MC_L1L2_L6D4),
.read_add_allproj(AP_L1L2_L6D4_MC_L1L2_L6D4_read_add),
.allprojin(AP_L1L2_L6D4_MC_L1L2_L6D4),
.read_add_allstub(AS_L6D4n4_MC_L1L2_L6D4_read_add),
.allstubin(AS_L6D4n4_MC_L1L2_L6D4),
.matchoutminus(MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus),
.matchoutplus(MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus),
.matchout1(MC_L1L2_L6D4_FM_L1L2_L6D4),
.valid_matchminus(MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus_wr_en),
.valid_match(MC_L1L2_L6D4_FM_L1L2_L6D4_wr_en),
.start(start8_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchTransceiver  MT_L3L4_Minus(
.number_in1(FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus_number),
.read_add1(FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus_read_add),
.proj1in(FM_L3L4_L1D3_ToMinus_MT_L3L4_Minus),
.number_in2(FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus_number),
.read_add2(FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus_read_add),
.proj2in(FM_L3L4_L1D4_ToMinus_MT_L3L4_Minus),
.number_in3(FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus_number),
.read_add3(FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus_read_add),
.proj3in(FM_L3L4_L2D3_ToMinus_MT_L3L4_Minus),
.number_in4(FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus_number),
.read_add4(FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus_read_add),
.proj4in(FM_L3L4_L2D4_ToMinus_MT_L3L4_Minus),
.number_in5(FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus_number),
.read_add5(FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus_read_add),
.proj5in(FM_L3L4_L5D3_ToMinus_MT_L3L4_Minus),
.number_in6(FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus_number),
.read_add6(FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus_read_add),
.proj6in(FM_L3L4_L5D4_ToMinus_MT_L3L4_Minus),
.number_in7(FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus_number),
.read_add7(FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus_read_add),
.proj7in(FM_L3L4_L6D3_ToMinus_MT_L3L4_Minus),
.number_in8(FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus_number),
.read_add8(FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus_read_add),
.proj8in(FM_L3L4_L6D4_ToMinus_MT_L3L4_Minus),
.valid_incomming_match_data_stream(MT_L3L4_Minus_From_DataStream_en),
.incomming_match_data_stream(MT_L3L4_Minus_From_DataStream),
.matchout1(MT_L3L4_Minus_FM_L3L4_L1_FromMinus),
.matchout2(MT_L3L4_Minus_FM_L3L4_L2_FromMinus),
.matchout3(MT_L3L4_Minus_FM_L3L4_L5_FromMinus),
.matchout4(MT_L3L4_Minus_FM_L3L4_L6_FromMinus),
.valid_matchout1(MT_L3L4_Minus_FM_L3L4_L1_FromMinus_wr_en),
.valid_matchout2(MT_L3L4_Minus_FM_L3L4_L2_FromMinus_wr_en),
.valid_matchout3(MT_L3L4_Minus_FM_L3L4_L5_FromMinus_wr_en),
.valid_matchout4(MT_L3L4_Minus_FM_L3L4_L6_FromMinus_wr_en),
.valid_match_data_stream(MT_L3L4_Minus_To_DataStream_en),
.match_data_stream(MT_L3L4_Minus_To_DataStream),
.start(start9_5),
.done(done9_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchTransceiver  MT_L5L6_Minus(
.number_in1(FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus_number),
.read_add1(FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus_read_add),
.proj1in(FM_L5L6_L1D3_ToMinus_MT_L5L6_Minus),
.number_in2(FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus_number),
.read_add2(FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus_read_add),
.proj2in(FM_L5L6_L1D4_ToMinus_MT_L5L6_Minus),
.number_in3(FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus_number),
.read_add3(FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus_read_add),
.proj3in(FM_L5L6_L2D3_ToMinus_MT_L5L6_Minus),
.number_in4(FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus_number),
.read_add4(FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus_read_add),
.proj4in(FM_L5L6_L2D4_ToMinus_MT_L5L6_Minus),
.number_in5(FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus_number),
.read_add5(FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus_read_add),
.proj5in(FM_L5L6_L3D3_ToMinus_MT_L5L6_Minus),
.number_in6(FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus_number),
.read_add6(FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus_read_add),
.proj6in(FM_L5L6_L3D4_ToMinus_MT_L5L6_Minus),
.number_in7(FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus_number),
.read_add7(FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus_read_add),
.proj7in(FM_L5L6_L4D3_ToMinus_MT_L5L6_Minus),
.number_in8(FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus_number),
.read_add8(FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus_read_add),
.proj8in(FM_L5L6_L4D4_ToMinus_MT_L5L6_Minus),
.valid_incomming_match_data_stream(MT_L5L6_Minus_From_DataStream_en),
.incomming_match_data_stream(MT_L5L6_Minus_From_DataStream),
.matchout1(MT_L5L6_Minus_FM_L5L6_L1_FromMinus),
.matchout2(MT_L5L6_Minus_FM_L5L6_L2_FromMinus),
.matchout3(MT_L5L6_Minus_FM_L5L6_L3_FromMinus),
.matchout4(MT_L5L6_Minus_FM_L5L6_L4_FromMinus),
.valid_matchout1(MT_L5L6_Minus_FM_L5L6_L1_FromMinus_wr_en),
.valid_matchout2(MT_L5L6_Minus_FM_L5L6_L2_FromMinus_wr_en),
.valid_matchout3(MT_L5L6_Minus_FM_L5L6_L3_FromMinus_wr_en),
.valid_matchout4(MT_L5L6_Minus_FM_L5L6_L4_FromMinus_wr_en),
.valid_match_data_stream(MT_L5L6_Minus_To_DataStream_en),
.match_data_stream(MT_L5L6_Minus_To_DataStream),
.start(start9_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchTransceiver  MT_L1L2_Minus(
.number_in1(FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus_number),
.read_add1(FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus_read_add),
.proj1in(FM_L1L2_L3D3_ToMinus_MT_L1L2_Minus),
.number_in2(FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus_number),
.read_add2(FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus_read_add),
.proj2in(FM_L1L2_L3D4_ToMinus_MT_L1L2_Minus),
.number_in3(FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus_number),
.read_add3(FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus_read_add),
.proj3in(FM_L1L2_L4D3_ToMinus_MT_L1L2_Minus),
.number_in4(FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus_number),
.read_add4(FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus_read_add),
.proj4in(FM_L1L2_L4D4_ToMinus_MT_L1L2_Minus),
.number_in5(FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus_number),
.read_add5(FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus_read_add),
.proj5in(FM_L1L2_L5D3_ToMinus_MT_L1L2_Minus),
.number_in6(FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus_number),
.read_add6(FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus_read_add),
.proj6in(FM_L1L2_L5D4_ToMinus_MT_L1L2_Minus),
.number_in7(FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus_number),
.read_add7(FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus_read_add),
.proj7in(FM_L1L2_L6D3_ToMinus_MT_L1L2_Minus),
.number_in8(FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus_number),
.read_add8(FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus_read_add),
.proj8in(FM_L1L2_L6D4_ToMinus_MT_L1L2_Minus),
.valid_incomming_match_data_stream(MT_L1L2_Minus_From_DataStream_en),
.incomming_match_data_stream(MT_L1L2_Minus_From_DataStream),
.matchout1(MT_L1L2_Minus_FM_L1L2_L3_FromMinus),
.matchout2(MT_L1L2_Minus_FM_L1L2_L4_FromMinus),
.matchout3(MT_L1L2_Minus_FM_L1L2_L5_FromMinus),
.matchout4(MT_L1L2_Minus_FM_L1L2_L6_FromMinus),
.valid_matchout1(MT_L1L2_Minus_FM_L1L2_L3_FromMinus_wr_en),
.valid_matchout2(MT_L1L2_Minus_FM_L1L2_L4_FromMinus_wr_en),
.valid_matchout3(MT_L1L2_Minus_FM_L1L2_L5_FromMinus_wr_en),
.valid_matchout4(MT_L1L2_Minus_FM_L1L2_L6_FromMinus_wr_en),
.valid_match_data_stream(MT_L1L2_Minus_To_DataStream_en),
.match_data_stream(MT_L1L2_Minus_To_DataStream),
.start(start9_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchTransceiver  MT_L3L4_Plus(
.number_in1(FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus_number),
.read_add1(FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus_read_add),
.proj1in(FM_L3L4_L1D3_ToPlus_MT_L3L4_Plus),
.number_in2(FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus_number),
.read_add2(FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus_read_add),
.proj2in(FM_L3L4_L1D4_ToPlus_MT_L3L4_Plus),
.number_in3(FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus_number),
.read_add3(FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus_read_add),
.proj3in(FM_L3L4_L2D3_ToPlus_MT_L3L4_Plus),
.number_in4(FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus_number),
.read_add4(FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus_read_add),
.proj4in(FM_L3L4_L2D4_ToPlus_MT_L3L4_Plus),
.number_in5(FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus_number),
.read_add5(FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus_read_add),
.proj5in(FM_L3L4_L5D3_ToPlus_MT_L3L4_Plus),
.number_in6(FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus_number),
.read_add6(FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus_read_add),
.proj6in(FM_L3L4_L5D4_ToPlus_MT_L3L4_Plus),
.number_in7(FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus_number),
.read_add7(FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus_read_add),
.proj7in(FM_L3L4_L6D3_ToPlus_MT_L3L4_Plus),
.number_in8(FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus_number),
.read_add8(FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus_read_add),
.proj8in(FM_L3L4_L6D4_ToPlus_MT_L3L4_Plus),
.valid_incomming_match_data_stream(MT_L3L4_Plus_From_DataStream_en),
.incomming_match_data_stream(MT_L3L4_Plus_From_DataStream),
.matchout1(MT_L3L4_Plus_FM_L3L4_L1_FromPlus),
.matchout2(MT_L3L4_Plus_FM_L3L4_L2_FromPlus),
.matchout3(MT_L3L4_Plus_FM_L3L4_L5_FromPlus),
.matchout4(MT_L3L4_Plus_FM_L3L4_L6_FromPlus),
.valid_matchout1(MT_L3L4_Plus_FM_L3L4_L1_FromPlus_wr_en),
.valid_matchout2(MT_L3L4_Plus_FM_L3L4_L2_FromPlus_wr_en),
.valid_matchout3(MT_L3L4_Plus_FM_L3L4_L5_FromPlus_wr_en),
.valid_matchout4(MT_L3L4_Plus_FM_L3L4_L6_FromPlus_wr_en),
.valid_match_data_stream(MT_L3L4_Plus_To_DataStream_en),
.match_data_stream(MT_L3L4_Plus_To_DataStream),
.start(start9_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchTransceiver  MT_L5L6_Plus(
.number_in1(FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus_number),
.read_add1(FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus_read_add),
.proj1in(FM_L5L6_L1D3_ToPlus_MT_L5L6_Plus),
.number_in2(FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus_number),
.read_add2(FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus_read_add),
.proj2in(FM_L5L6_L1D4_ToPlus_MT_L5L6_Plus),
.number_in3(FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus_number),
.read_add3(FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus_read_add),
.proj3in(FM_L5L6_L2D3_ToPlus_MT_L5L6_Plus),
.number_in4(FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus_number),
.read_add4(FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus_read_add),
.proj4in(FM_L5L6_L2D4_ToPlus_MT_L5L6_Plus),
.number_in5(FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus_number),
.read_add5(FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus_read_add),
.proj5in(FM_L5L6_L3D3_ToPlus_MT_L5L6_Plus),
.number_in6(FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus_number),
.read_add6(FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus_read_add),
.proj6in(FM_L5L6_L3D4_ToPlus_MT_L5L6_Plus),
.number_in7(FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus_number),
.read_add7(FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus_read_add),
.proj7in(FM_L5L6_L4D3_ToPlus_MT_L5L6_Plus),
.number_in8(FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus_number),
.read_add8(FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus_read_add),
.proj8in(FM_L5L6_L4D4_ToPlus_MT_L5L6_Plus),
.valid_incomming_match_data_stream(MT_L5L6_Plus_From_DataStream_en),
.incomming_match_data_stream(MT_L5L6_Plus_From_DataStream),
.matchout1(MT_L5L6_Plus_FM_L5L6_L1_FromPlus),
.matchout2(MT_L5L6_Plus_FM_L5L6_L2_FromPlus),
.matchout3(MT_L5L6_Plus_FM_L5L6_L3_FromPlus),
.matchout4(MT_L5L6_Plus_FM_L5L6_L4_FromPlus),
.valid_matchout1(MT_L5L6_Plus_FM_L5L6_L1_FromPlus_wr_en),
.valid_matchout2(MT_L5L6_Plus_FM_L5L6_L2_FromPlus_wr_en),
.valid_matchout3(MT_L5L6_Plus_FM_L5L6_L3_FromPlus_wr_en),
.valid_matchout4(MT_L5L6_Plus_FM_L5L6_L4_FromPlus_wr_en),
.valid_match_data_stream(MT_L5L6_Plus_To_DataStream_en),
.match_data_stream(MT_L5L6_Plus_To_DataStream),
.start(start9_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


MatchTransceiver  MT_L1L2_Plus(
.number_in1(FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus_number),
.read_add1(FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus_read_add),
.proj1in(FM_L1L2_L3D3_ToPlus_MT_L1L2_Plus),
.number_in2(FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus_number),
.read_add2(FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus_read_add),
.proj2in(FM_L1L2_L3D4_ToPlus_MT_L1L2_Plus),
.number_in3(FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus_number),
.read_add3(FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus_read_add),
.proj3in(FM_L1L2_L4D3_ToPlus_MT_L1L2_Plus),
.number_in4(FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus_number),
.read_add4(FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus_read_add),
.proj4in(FM_L1L2_L4D4_ToPlus_MT_L1L2_Plus),
.number_in5(FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus_number),
.read_add5(FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus_read_add),
.proj5in(FM_L1L2_L5D3_ToPlus_MT_L1L2_Plus),
.number_in6(FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus_number),
.read_add6(FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus_read_add),
.proj6in(FM_L1L2_L5D4_ToPlus_MT_L1L2_Plus),
.number_in7(FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus_number),
.read_add7(FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus_read_add),
.proj7in(FM_L1L2_L6D3_ToPlus_MT_L1L2_Plus),
.number_in8(FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus_number),
.read_add8(FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus_read_add),
.proj8in(FM_L1L2_L6D4_ToPlus_MT_L1L2_Plus),
.valid_incomming_match_data_stream(MT_L1L2_Plus_From_DataStream_en),
.incomming_match_data_stream(MT_L1L2_Plus_From_DataStream),
.matchout1(MT_L1L2_Plus_FM_L1L2_L3_FromPlus),
.matchout2(MT_L1L2_Plus_FM_L1L2_L4_FromPlus),
.matchout3(MT_L1L2_Plus_FM_L1L2_L5_FromPlus),
.matchout4(MT_L1L2_Plus_FM_L1L2_L6_FromPlus),
.valid_matchout1(MT_L1L2_Plus_FM_L1L2_L3_FromPlus_wr_en),
.valid_matchout2(MT_L1L2_Plus_FM_L1L2_L4_FromPlus_wr_en),
.valid_matchout3(MT_L1L2_Plus_FM_L1L2_L5_FromPlus_wr_en),
.valid_matchout4(MT_L1L2_Plus_FM_L1L2_L6_FromPlus_wr_en),
.valid_match_data_stream(MT_L1L2_Plus_To_DataStream_en),
.match_data_stream(MT_L1L2_Plus_To_DataStream),
.start(start9_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


FitTrack  FT_L1L2(
.number1in1(FM_L1L2_L3D3_FT_L1L2_number),
.read_add1in1(FM_L1L2_L3D3_FT_L1L2_read_add),
.read_en1in1(FM_L1L2_L3D3_FT_L1L2_read_en),
.fullmatch1in1(FM_L1L2_L3D3_FT_L1L2),
.number1in2(FM_L1L2_L3D4_FT_L1L2_number),
.read_add1in2(FM_L1L2_L3D4_FT_L1L2_read_add),
.read_en1in2(FM_L1L2_L3D4_FT_L1L2_read_en),
.fullmatch1in2(FM_L1L2_L3D4_FT_L1L2),
.number2in1(FM_L1L2_L4D3_FT_L1L2_number),
.read_add2in1(FM_L1L2_L4D3_FT_L1L2_read_add),
.read_en2in1(FM_L1L2_L4D3_FT_L1L2_read_en),
.fullmatch2in1(FM_L1L2_L4D3_FT_L1L2),
.number2in2(FM_L1L2_L4D4_FT_L1L2_number),
.read_add2in2(FM_L1L2_L4D4_FT_L1L2_read_add),
.read_en2in2(FM_L1L2_L4D4_FT_L1L2_read_en),
.fullmatch2in2(FM_L1L2_L4D4_FT_L1L2),
.number3in1(FM_L1L2_L5D3_FT_L1L2_number),
.read_add3in1(FM_L1L2_L5D3_FT_L1L2_read_add),
.read_en3in1(FM_L1L2_L5D3_FT_L1L2_read_en),
.fullmatch3in1(FM_L1L2_L5D3_FT_L1L2),
.number3in2(FM_L1L2_L5D4_FT_L1L2_number),
.read_add3in2(FM_L1L2_L5D4_FT_L1L2_read_add),
.read_en3in2(FM_L1L2_L5D4_FT_L1L2_read_en),
.fullmatch3in2(FM_L1L2_L5D4_FT_L1L2),
.number4in1(FM_L1L2_L6D3_FT_L1L2_number),
.read_add4in1(FM_L1L2_L6D3_FT_L1L2_read_add),
.read_en4in1(FM_L1L2_L6D3_FT_L1L2_read_en),
.fullmatch4in1(FM_L1L2_L6D3_FT_L1L2),
.number4in2(FM_L1L2_L6D4_FT_L1L2_number),
.read_add4in2(FM_L1L2_L6D4_FT_L1L2_read_add),
.read_en4in2(FM_L1L2_L6D4_FT_L1L2_read_en),
.fullmatch4in2(FM_L1L2_L6D4_FT_L1L2),
.number1in3(FM_L1L2_L3_FromPlus_FT_L1L2_number),
.read_add1in3(FM_L1L2_L3_FromPlus_FT_L1L2_read_add),
.read_en1in3(FM_L1L2_L3_FromPlus_FT_L1L2_read_en),
.fullmatch1in3(FM_L1L2_L3_FromPlus_FT_L1L2),
.number2in3(FM_L1L2_L4_FromPlus_FT_L1L2_number),
.read_add2in3(FM_L1L2_L4_FromPlus_FT_L1L2_read_add),
.read_en2in3(FM_L1L2_L4_FromPlus_FT_L1L2_read_en),
.fullmatch2in3(FM_L1L2_L4_FromPlus_FT_L1L2),
.number3in3(FM_L1L2_L5_FromPlus_FT_L1L2_number),
.read_add3in3(FM_L1L2_L5_FromPlus_FT_L1L2_read_add),
.read_en3in3(FM_L1L2_L5_FromPlus_FT_L1L2_read_en),
.fullmatch3in3(FM_L1L2_L5_FromPlus_FT_L1L2),
.number4in3(FM_L1L2_L6_FromPlus_FT_L1L2_number),
.read_add4in3(FM_L1L2_L6_FromPlus_FT_L1L2_read_add),
.read_en4in3(FM_L1L2_L6_FromPlus_FT_L1L2_read_en),
.fullmatch4in3(FM_L1L2_L6_FromPlus_FT_L1L2),
.number1in4(FM_L1L2_L3_FromMinus_FT_L1L2_number),
.read_add1in4(FM_L1L2_L3_FromMinus_FT_L1L2_read_add),
.read_en1in4(FM_L1L2_L3_FromMinus_FT_L1L2_read_en),
.fullmatch1in4(FM_L1L2_L3_FromMinus_FT_L1L2),
.number2in4(FM_L1L2_L4_FromMinus_FT_L1L2_number),
.read_add2in4(FM_L1L2_L4_FromMinus_FT_L1L2_read_add),
.read_en2in4(FM_L1L2_L4_FromMinus_FT_L1L2_read_en),
.fullmatch2in4(FM_L1L2_L4_FromMinus_FT_L1L2),
.number3in4(FM_L1L2_L5_FromMinus_FT_L1L2_number),
.read_add3in4(FM_L1L2_L5_FromMinus_FT_L1L2_read_add),
.read_en3in4(FM_L1L2_L5_FromMinus_FT_L1L2_read_en),
.fullmatch3in4(FM_L1L2_L5_FromMinus_FT_L1L2),
.number4in4(FM_L1L2_L6_FromMinus_FT_L1L2_number),
.read_add4in4(FM_L1L2_L6_FromMinus_FT_L1L2_read_add),
.read_en4in4(FM_L1L2_L6_FromMinus_FT_L1L2_read_en),
.fullmatch4in4(FM_L1L2_L6_FromMinus_FT_L1L2),
.read_add_pars1(TPAR_L1D3L2D3_FT_L1L2_read_add),
.tpar1in(TPAR_L1D3L2D3_FT_L1L2),
.read_add_pars2(TPAR_L1D4L2D4_FT_L1L2_read_add),
.tpar2in(TPAR_L1D4L2D4_FT_L1L2),
.read_add_pars3(TPAR_L1D3L2D4_FT_L1L2_read_add),
.tpar3in(TPAR_L1D3L2D4_FT_L1L2),
.trackout(FT_L1L2_TF_L1L2),
.valid_fit(FT_L1L2_TF_L1L2_wr_en),
.start(start10_5),
.done(done10_0),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


FitTrack  FT_L3L4(
.number1in1(FM_L3L4_L1D3_FT_L3L4_number),
.read_add1in1(FM_L3L4_L1D3_FT_L3L4_read_add),
.read_en1in1(FM_L3L4_L1D3_FT_L3L4_read_en),
.fullmatch1in1(FM_L3L4_L1D3_FT_L3L4),
.number1in2(FM_L3L4_L1D4_FT_L3L4_number),
.read_add1in2(FM_L3L4_L1D4_FT_L3L4_read_add),
.read_en1in2(FM_L3L4_L1D4_FT_L3L4_read_en),
.fullmatch1in2(FM_L3L4_L1D4_FT_L3L4),
.number2in1(FM_L3L4_L2D3_FT_L3L4_number),
.read_add2in1(FM_L3L4_L2D3_FT_L3L4_read_add),
.read_en2in1(FM_L3L4_L2D3_FT_L3L4_read_en),
.fullmatch2in1(FM_L3L4_L2D3_FT_L3L4),
.number2in2(FM_L3L4_L2D4_FT_L3L4_number),
.read_add2in2(FM_L3L4_L2D4_FT_L3L4_read_add),
.read_en2in2(FM_L3L4_L2D4_FT_L3L4_read_en),
.fullmatch2in2(FM_L3L4_L2D4_FT_L3L4),
.number3in1(FM_L3L4_L5D3_FT_L3L4_number),
.read_add3in1(FM_L3L4_L5D3_FT_L3L4_read_add),
.read_en3in1(FM_L3L4_L5D3_FT_L3L4_read_en),
.fullmatch3in1(FM_L3L4_L5D3_FT_L3L4),
.number3in2(FM_L3L4_L5D4_FT_L3L4_number),
.read_add3in2(FM_L3L4_L5D4_FT_L3L4_read_add),
.read_en3in2(FM_L3L4_L5D4_FT_L3L4_read_en),
.fullmatch3in2(FM_L3L4_L5D4_FT_L3L4),
.number4in1(FM_L3L4_L6D3_FT_L3L4_number),
.read_add4in1(FM_L3L4_L6D3_FT_L3L4_read_add),
.read_en4in1(FM_L3L4_L6D3_FT_L3L4_read_en),
.fullmatch4in1(FM_L3L4_L6D3_FT_L3L4),
.number4in2(FM_L3L4_L6D4_FT_L3L4_number),
.read_add4in2(FM_L3L4_L6D4_FT_L3L4_read_add),
.read_en4in2(FM_L3L4_L6D4_FT_L3L4_read_en),
.fullmatch4in2(FM_L3L4_L6D4_FT_L3L4),
.number1in3(FM_L3L4_L1_FromMinus_FT_L3L4_number),
.read_add1in3(FM_L3L4_L1_FromMinus_FT_L3L4_read_add),
.read_en1in3(FM_L3L4_L1_FromMinus_FT_L3L4_read_en),
.fullmatch1in3(FM_L3L4_L1_FromMinus_FT_L3L4),
.number2in3(FM_L3L4_L2_FromMinus_FT_L3L4_number),
.read_add2in3(FM_L3L4_L2_FromMinus_FT_L3L4_read_add),
.read_en2in3(FM_L3L4_L2_FromMinus_FT_L3L4_read_en),
.fullmatch2in3(FM_L3L4_L2_FromMinus_FT_L3L4),
.number3in3(FM_L3L4_L5_FromMinus_FT_L3L4_number),
.read_add3in3(FM_L3L4_L5_FromMinus_FT_L3L4_read_add),
.read_en3in3(FM_L3L4_L5_FromMinus_FT_L3L4_read_en),
.fullmatch3in3(FM_L3L4_L5_FromMinus_FT_L3L4),
.number4in3(FM_L3L4_L6_FromMinus_FT_L3L4_number),
.read_add4in3(FM_L3L4_L6_FromMinus_FT_L3L4_read_add),
.read_en4in3(FM_L3L4_L6_FromMinus_FT_L3L4_read_en),
.fullmatch4in3(FM_L3L4_L6_FromMinus_FT_L3L4),
.number1in4(FM_L3L4_L1_FromPlus_FT_L3L4_number),
.read_add1in4(FM_L3L4_L1_FromPlus_FT_L3L4_read_add),
.read_en1in4(FM_L3L4_L1_FromPlus_FT_L3L4_read_en),
.fullmatch1in4(FM_L3L4_L1_FromPlus_FT_L3L4),
.number2in4(FM_L3L4_L2_FromPlus_FT_L3L4_number),
.read_add2in4(FM_L3L4_L2_FromPlus_FT_L3L4_read_add),
.read_en2in4(FM_L3L4_L2_FromPlus_FT_L3L4_read_en),
.fullmatch2in4(FM_L3L4_L2_FromPlus_FT_L3L4),
.number3in4(FM_L3L4_L5_FromPlus_FT_L3L4_number),
.read_add3in4(FM_L3L4_L5_FromPlus_FT_L3L4_read_add),
.read_en3in4(FM_L3L4_L5_FromPlus_FT_L3L4_read_en),
.fullmatch3in4(FM_L3L4_L5_FromPlus_FT_L3L4),
.number4in4(FM_L3L4_L6_FromPlus_FT_L3L4_number),
.read_add4in4(FM_L3L4_L6_FromPlus_FT_L3L4_read_add),
.read_en4in4(FM_L3L4_L6_FromPlus_FT_L3L4_read_en),
.fullmatch4in4(FM_L3L4_L6_FromPlus_FT_L3L4),
.read_add_pars1(TPAR_L3D3L4D3_FT_L3L4_read_add),
.tpar1in(TPAR_L3D3L4D3_FT_L3L4),
.read_add_pars2(TPAR_L3D3L4D4_FT_L3L4_read_add),
.tpar2in(TPAR_L3D3L4D4_FT_L3L4),
.read_add_pars3(TPAR_L3D4L4D4_FT_L3L4_read_add),
.tpar3in(TPAR_L3D4L4D4_FT_L3L4),
.trackout(FT_L3L4_TF_L3L4),
.valid_fit(FT_L3L4_TF_L3L4_wr_en),
.start(start10_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);


FitTrack  FT_L5L6(
.number1in1(FM_L5L6_L1D3_FT_L5L6_number),
.read_add1in1(FM_L5L6_L1D3_FT_L5L6_read_add),
.read_en1in1(FM_L5L6_L1D3_FT_L5L6_read_en),
.fullmatch1in1(FM_L5L6_L1D3_FT_L5L6),
.number1in2(FM_L5L6_L1D4_FT_L5L6_number),
.read_add1in2(FM_L5L6_L1D4_FT_L5L6_read_add),
.read_en1in2(FM_L5L6_L1D4_FT_L5L6_read_en),
.fullmatch1in2(FM_L5L6_L1D4_FT_L5L6),
.number2in1(FM_L5L6_L2D3_FT_L5L6_number),
.read_add2in1(FM_L5L6_L2D3_FT_L5L6_read_add),
.read_en2in1(FM_L5L6_L2D3_FT_L5L6_read_en),
.fullmatch2in1(FM_L5L6_L2D3_FT_L5L6),
.number2in2(FM_L5L6_L2D4_FT_L5L6_number),
.read_add2in2(FM_L5L6_L2D4_FT_L5L6_read_add),
.read_en2in2(FM_L5L6_L2D4_FT_L5L6_read_en),
.fullmatch2in2(FM_L5L6_L2D4_FT_L5L6),
.number3in1(FM_L5L6_L3D3_FT_L5L6_number),
.read_add3in1(FM_L5L6_L3D3_FT_L5L6_read_add),
.read_en3in1(FM_L5L6_L3D3_FT_L5L6_read_en),
.fullmatch3in1(FM_L5L6_L3D3_FT_L5L6),
.number3in2(FM_L5L6_L3D4_FT_L5L6_number),
.read_add3in2(FM_L5L6_L3D4_FT_L5L6_read_add),
.read_en3in2(FM_L5L6_L3D4_FT_L5L6_read_en),
.fullmatch3in2(FM_L5L6_L3D4_FT_L5L6),
.number4in1(FM_L5L6_L4D3_FT_L5L6_number),
.read_add4in1(FM_L5L6_L4D3_FT_L5L6_read_add),
.read_en4in1(FM_L5L6_L4D3_FT_L5L6_read_en),
.fullmatch4in1(FM_L5L6_L4D3_FT_L5L6),
.number4in2(FM_L5L6_L4D4_FT_L5L6_number),
.read_add4in2(FM_L5L6_L4D4_FT_L5L6_read_add),
.read_en4in2(FM_L5L6_L4D4_FT_L5L6_read_en),
.fullmatch4in2(FM_L5L6_L4D4_FT_L5L6),
.number1in3(FM_L5L6_L1_FromPlus_FT_L5L6_number),
.read_add1in3(FM_L5L6_L1_FromPlus_FT_L5L6_read_add),
.read_en1in3(FM_L5L6_L1_FromPlus_FT_L5L6_read_en),
.fullmatch1in3(FM_L5L6_L1_FromPlus_FT_L5L6),
.number2in3(FM_L5L6_L2_FromPlus_FT_L5L6_number),
.read_add2in3(FM_L5L6_L2_FromPlus_FT_L5L6_read_add),
.read_en2in3(FM_L5L6_L2_FromPlus_FT_L5L6_read_en),
.fullmatch2in3(FM_L5L6_L2_FromPlus_FT_L5L6),
.number3in3(FM_L5L6_L3_FromPlus_FT_L5L6_number),
.read_add3in3(FM_L5L6_L3_FromPlus_FT_L5L6_read_add),
.read_en3in3(FM_L5L6_L3_FromPlus_FT_L5L6_read_en),
.fullmatch3in3(FM_L5L6_L3_FromPlus_FT_L5L6),
.number4in3(FM_L5L6_L4_FromPlus_FT_L5L6_number),
.read_add4in3(FM_L5L6_L4_FromPlus_FT_L5L6_read_add),
.read_en4in3(FM_L5L6_L4_FromPlus_FT_L5L6_read_en),
.fullmatch4in3(FM_L5L6_L4_FromPlus_FT_L5L6),
.number1in4(FM_L5L6_L1_FromMinus_FT_L5L6_number),
.read_add1in4(FM_L5L6_L1_FromMinus_FT_L5L6_read_add),
.read_en1in4(FM_L5L6_L1_FromMinus_FT_L5L6_read_en),
.fullmatch1in4(FM_L5L6_L1_FromMinus_FT_L5L6),
.number2in4(FM_L5L6_L2_FromMinus_FT_L5L6_number),
.read_add2in4(FM_L5L6_L2_FromMinus_FT_L5L6_read_add),
.read_en2in4(FM_L5L6_L2_FromMinus_FT_L5L6_read_en),
.fullmatch2in4(FM_L5L6_L2_FromMinus_FT_L5L6),
.number3in4(FM_L5L6_L3_FromMinus_FT_L5L6_number),
.read_add3in4(FM_L5L6_L3_FromMinus_FT_L5L6_read_add),
.read_en3in4(FM_L5L6_L3_FromMinus_FT_L5L6_read_en),
.fullmatch3in4(FM_L5L6_L3_FromMinus_FT_L5L6),
.number4in4(FM_L5L6_L4_FromMinus_FT_L5L6_number),
.read_add4in4(FM_L5L6_L4_FromMinus_FT_L5L6_read_add),
.read_en4in4(FM_L5L6_L4_FromMinus_FT_L5L6_read_en),
.fullmatch4in4(FM_L5L6_L4_FromMinus_FT_L5L6),
.read_add_pars1(TPAR_L5D3L6D3_FT_L5L6_read_add),
.tpar1in(TPAR_L5D3L6D3_FT_L5L6),
.read_add_pars2(TPAR_L5D4L6D4_FT_L5L6_read_add),
.tpar2in(TPAR_L5D4L6D4_FT_L5L6),
.read_add_pars3(TPAR_L5D3L6D4_FT_L5L6_read_add),
.tpar3in(TPAR_L5D3L6D4_FT_L5L6),
.trackout(FT_L5L6_TF_L5L6),
.valid_fit(FT_L5L6_TF_L5L6_wr_en),
.start(start10_5),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [31:0] reader_out;

//reader reader1(

//.read_add1(TPAR_L1D3L2D3_FT_L1L2_read_add),
//.read_add2(TPROJ_L1D3L2D3_L3_PR_L3D3_L1L2_read_add),
//.read_add3(SL1_L3D3_VMR_L3D3_read_add),
//.read_add4(SL1_L4D3_VMR_L4D3_read_add),
//.read_add5(SL1_L5D3_VMR_L5D3_read_add),

//.number_in1(TPAR_L1D3L2D3_FT_L1L2_number),
//.number_in2(TPROJ_L1D3L2D3_L3_PR_L3D3_L1L2_number),
//.number_in3(SL1_L3D3_VMR_L3D3_number),
//.number_in4(SL1_L4D3_VMR_L4D3_number),
//.number_in5(SL1_L5D3_VMR_L5D3_number),

//.input1(TPAR_L1D3L2D3_FT_L1L2),
//.input2(TPROJ_L1D3L2D3_L3_PR_L3D3_L1L2),
//.input3(SL1_L3D3_VMR_L3D3),
//.input4(SL1_L4D3_VMR_L4D3),
//.input5(SL1_L5D3_VMR_L5D3),

//.clk(clk),
//.reset(reset),
//.en_proc(enable_gen),
//.io_clk(io_clk),
//.io_sel(io_sel_R3_io_block),
//.io_addr(io_addr[15:0]),
//.io_sync(io_sync),
//.io_rd_en(io_rd_en),
//.io_wr_en(io_wr_en),
//.io_wr_data(io_wr_data[31:0]),
//.io_rd_data(reader_out),
//.io_rd_ack(reader_ack),
//.BX(BX[2:0]),
//.first_clk(first_clk),
//.not_first_clk(not_first_clk)
//);

wire InputLink_R1Link1_io_rd_ack , InputLink_R1Link2_io_rd_ack , InputLink_R1Link3_io_rd_ack;
wire TPars_L1L2_io_rd_ack , TPars_L3L4_io_rd_ack , TPars_L5L6_io_rd_ack;
// readback mux
// If a particular block is addressed, connect that block's signals
// to the 'rdbk' output. At the same time, assert 'rdbk_sel' to tell downstream muxes to
// use the 'rdbk' from this module as their source of data.
reg [31:0] io_rd_data_reg;
assign io_rd_data = io_rd_data_reg;
// Assert 'io_rd_ack' if any module is asserting its 'rd_ack'.
reg io_rd_ack_reg;
assign io_rd_ack = io_rd_ack_reg;
always @ (posedge io_clk) begin
io_rd_ack_reg <= InputLink_R1Link1_io_rd_ack | InputLink_R1Link2_io_rd_ack | InputLink_R1Link3_io_rd_ack |
TPars_L1L2_io_rd_ack | TPars_L3L4_io_rd_ack | TPars_L5L6_io_rd_ack;
end
// Route the selected register to the 'rdbk' output.
always @(posedge io_clk) begin
if (InputLink_R1Link1_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link1_io_rd_data[31:0];
if (InputLink_R1Link2_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link2_io_rd_data[31:0];
if (InputLink_R1Link3_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link3_io_rd_data[31:0];
if (TPars_L1L2_io_sel) io_rd_data_reg[31:0] <= TPars_L1L2_io_rd_data[31:0];
if (TPars_L3L4_io_sel) io_rd_data_reg[31:0] <= TPars_L3L4_io_rd_data[31:0];
if (TPars_L5L6_io_sel) io_rd_data_reg[31:0] <= TPars_L5L6_io_rd_data[31:0];
//if (reader_ack)    io_rd_data_reg <= reader_out;
end

endmodule

