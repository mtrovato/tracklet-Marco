`timescale 1ns / 1ps
`include "constants.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/28/2014 03:18:24 PM
// Design Name: 
// Module Name: VMStubs
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module VMStubs(
    input clk,
    input reset,
    input en_proc,
    input [1:0] start,
    output [1:0] done,
    
    input [18:0] data_in,
    input enable,
    
    output [5:0] number_out,
    input [4+`MEM_SIZE:0] read_add,
    output reg [18:0] data_out
    );

    parameter engine="Tracklet";

    reg [18:0] data_in_dly;
    reg [`MEM_SIZE:0] wr_add;
    reg wr_en;
    
    reg [4:0] BX_pipe;
    reg [4:0] BX_dly;
    reg first_clk_pipe;
    
    reg [1:0] rst_pipe;
    
    initial begin
        BX_pipe = 5'b11111;
    end
    
    always @(posedge clk) begin
        rst_pipe <= start;     // use the top bit of start as pipelined reset
        BX_dly <= BX_pipe;    
        if(rst_pipe[1])
            BX_pipe <= 5'b11111; 
        else begin
            if(rst_pipe[0]) begin
                BX_pipe <= BX_pipe + 1'b1;
                first_clk_pipe <= 1'b1;
            end
            else begin
                first_clk_pipe <= 1'b0;
            end
        end
    end
    
    wire [18:0] pre_data_out;
    
    always @(posedge clk) begin
        data_in_dly <= data_in;
        if(first_clk_pipe) begin
            wr_add <= {`MEM_SIZE+1{1'b1}};
            //number_out <= wr_add + 1'b1;
        end
        else begin
            if(enable & data_in[15:10] < 6'b011111) begin
                wr_add <= wr_add + 1'b1;
                wr_en <= 1'b1;
            end
            else begin
                wr_add <= wr_add;
                wr_en <= 1'b0;
            end
        end
        data_out <= pre_data_out;
    end
    
    pipe_delay #(.STAGES(`tmux+2), .WIDTH(3))
               done_delay(.pipe_in(), .pipe_out(), .clk(clk),
               .val_in(start), .val_out(done));
   // Could make this a DRAM for Tracklet Engines
   
   generate
       if(engine=="Match")
           Memory #(
               .RAM_WIDTH(19),                       // Specify RAM data width
               .RAM_DEPTH(2**(`MEM_SIZE+5)),                     // Specify RAM depth (number of entries)
               .RAM_PERFORMANCE("HIGH_PERFORMANCE"), // Select "HIGH_PERFORMANCE" or "LOW_LATENCY" 
               .INIT_FILE("")                        // Specify name/location of RAM initialization file if using one (leave blank if not)
             ) VMStubME (
               .addra({BX_dly[4:0],wr_add[`MEM_SIZE-1:0]}),    // Write address bus, width determined from RAM_DEPTH
               .addrb(read_add[(`MEM_SIZE+5)-1:0]),    // Read address bus, width determined from RAM_DEPTH
               .dina(data_in_dly),      // RAM input data, width determined from RAM_WIDTH
               .clka(clk),      // Write clock
               .clkb(clk),      // Read clock
               .wea(wr_en),        // Write enable
               .enb(1'b1),        // Read Enable, for additional power savings, disable when not in use
               .rstb(rst_pipe),      // Output reset (does not affect memory contents)
               .regceb(1'b1),  // Output register enable
               .doutb(pre_data_out)     // RAM output data, width determined from RAM_WIDTH
               );
       else
           reg_array #(
             //Memory #(
                 .RAM_WIDTH(19),                       // Specify RAM data width
                 .RAM_DEPTH(2**(`MEM_SIZE+1)),                     // Specify RAM depth (number of entries)
                 .INIT_FILE("") //"full.txt")                        // Specify name/location of RAM initialization file if using one (leave blank if not)
               ) VMStubTE (
                 .addra({BX_dly[0],wr_add[`MEM_SIZE-1:0]}),    // Write address bus, width determined from RAM_DEPTH
                 .addrb(read_add[`MEM_SIZE:0]),    // Read address bus, width determined from RAM_DEPTH
                 .dina(data_in_dly),      // RAM input data, width determined from RAM_WIDTH
                 .clka(clk),      // Write clock
                 .clkb(clk),      // Read clock
                 .wea(wr_en),        // Write enable
                 //.enb(1'b1),        // Read Enable, for additional power savings, disable when not in use // Maybe don't read add = 6'h3f?
                 .rstb(rst_pipe),      // Output reset (does not affect memory contents)
                 .regceb(1'b1),  // Output register enable
                 //.doutb(pre_data_out)     // RAM output data, width determined from RAM_WIDTH
                 .doutb(pre_data_out)
             );
   endgenerate
    
        
    reg_array #(
      //Memory #(
              .RAM_WIDTH(6),                       // Specify RAM data width
              .RAM_DEPTH(32),                     // Specify RAM depth (number of entries)
              .INIT_FILE("") //"full.txt")                        // Specify name/location of RAM initialization file if using one (leave blank if not)
            ) Number_out (
              .addra(BX_dly),    // Write address bus, width determined from RAM_DEPTH
              .addrb(read_add[9:5]),    // Read address bus, width determined from RAM_DEPTH
              .dina(wr_add+1'b1),      // RAM input data, width determined from RAM_WIDTH
              .clka(clk),      // Write clock
              .clkb(clk),      // Read clock
              .wea(1'b1),        // Write enable
              //.enb(1'b1),        // Read Enable, for additional power savings, disable when not in use // Maybe don't read add = 6'h3f?
              .rstb(rst_pipe),      // Output reset (does not affect memory contents)
              .regceb(1'b1),  // Output register enable
              //.doutb(pre_data_out)     // RAM output data, width determined from RAM_WIDTH
              .doutb(number_out)
      );
    
endmodule
