
`timescale 1ns / 1ps
`include "constants.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 09/28/2014 11:01:39 AM
// Design Name:
// Module Name: Tracklet_processing
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module Tracklet_processingD3D4(
input clk,
input clk_new, //MT			   
input reset,
input en_proc,
// programming interface
// inputs
input wire io_clk,                    // programming clock
input wire io_sel,                    // this module has been selected for an I/O operation
input wire io_sync,
// start the I/O operation
input wire [15:0] io_addr,        // slave address, memory or register. Top 12 bits already consumed.
input wire io_rd_en,                // this is a read operation
input wire io_wr_en,                // this is a write operation
input wire [31:0] io_wr_data,    // data to write for write operations
// outputs
output wire [31:0] io_rd_data,    // data returned for read operations
output wire io_rd_ack,                // 'read' data from this module is ready
//clocks
input wire [2:0] BX,
input wire first_clk,
input wire not_first_clk,
// inputs
input [31:0] input_link1_reg1,
input [31:0] input_link1_reg2,
input [31:0] input_link2_reg1,
input [31:0] input_link2_reg2,
input [31:0] input_link3_reg1,
input [31:0] input_link3_reg2,
input [31:0] input_link4_reg1,
input [31:0] input_link4_reg2,
input [31:0] input_link5_reg1,
input [31:0] input_link5_reg2,
input [31:0] input_link6_reg1,
input [31:0] input_link6_reg2,
input [31:0] input_link7_reg1,
input [31:0] input_link7_reg2,
input [31:0] input_link8_reg1,
input [31:0] input_link8_reg2,
input [31:0] input_link9_reg1,
input [31:0] input_link9_reg2,
// outputs
input [15:0] BRAM_OUTPUT_addr, // 1 for now, add more later
input BRAM_OUTPUT_clk,
input [31:0] BRAM_OUTPUT_din,
output [31:0] BRAM_OUTPUT_dout,
input BRAM_OUTPUT_en,
input BRAM_OUTPUT_rst,
input [3:0] BRAM_OUTPUT_we,
// Projections L3F3F5
output wire [54:0] PT_L3F3F5_Plus_To_DataStream,
output wire PT_L3F3F5_Plus_To_DataStream_en,
output wire [54:0] PT_L3F3F5_Minus_To_DataStream,
output wire PT_L3F3F5_Minus_To_DataStream_en,
input wire [54:0] PT_L3F3F5_Plus_From_DataStream,
input wire PT_L3F3F5_Plus_From_DataStream_en,
input wire [54:0] PT_L3F3F5_Minus_From_DataStream,
input wire PT_L3F3F5_Minus_From_DataStream_en,
// Projections L2L4F2
output wire [54:0] PT_L2L4F2_Plus_To_DataStream,
output wire PT_L2L4F2_Plus_To_DataStream_en,
output wire [54:0] PT_L2L4F2_Minus_To_DataStream,
output wire PT_L2L4F2_Minus_To_DataStream_en,
input wire [54:0] PT_L2L4F2_Plus_From_DataStream,
input wire PT_L2L4F2_Plus_From_DataStream_en,
input wire [54:0] PT_L2L4F2_Minus_From_DataStream,
input wire PT_L2L4F2_Minus_From_DataStream_en,
// Projections F1L5
output wire [54:0] PT_F1L5_Plus_To_DataStream,
output wire PT_F1L5_Plus_To_DataStream_en,
output wire [54:0] PT_F1L5_Minus_To_DataStream,
output wire PT_F1L5_Minus_To_DataStream_en,
input wire [54:0] PT_F1L5_Plus_From_DataStream,
input wire PT_F1L5_Plus_From_DataStream_en,
input wire [54:0] PT_F1L5_Minus_From_DataStream,
input wire PT_F1L5_Minus_From_DataStream_en,
// Projections L1L6F4
output wire [54:0] PT_L1L6F4_Plus_To_DataStream,
output wire PT_L1L6F4_Plus_To_DataStream_en,
output wire [54:0] PT_L1L6F4_Minus_To_DataStream,
output wire PT_L1L6F4_Minus_To_DataStream_en,
input wire [54:0] PT_L1L6F4_Plus_From_DataStream,
input wire PT_L1L6F4_Plus_From_DataStream_en,
input wire [54:0] PT_L1L6F4_Minus_From_DataStream,
input wire PT_L1L6F4_Minus_From_DataStream_en,
// Matches Disk
output wire [44:0] MT_FDSK_Minus_To_DataStream,
output wire MT_FDSK_Minus_To_DataStream_en,
output wire [44:0] MT_FDSK_Plus_To_DataStream,
output wire MT_FDSK_Plus_To_DataStream_en,
input wire [44:0] MT_FDSK_Plus_From_DataStream,
input wire MT_FDSK_Plus_From_DataStream_en,
input wire [44:0] MT_FDSK_Minus_From_DataStream,
input wire MT_FDSK_Minus_From_DataStream_en,
// Matches Layer
output wire [44:0] MT_Layr_Plus_To_DataStream,
output wire MT_Layr_Plus_To_DataStream_en,
output wire [44:0] MT_Layr_Minus_To_DataStream,
output wire MT_Layr_Minus_To_DataStream_en,
input wire [44:0] MT_Layr_Plus_From_DataStream,
input wire MT_Layr_Plus_From_DataStream_en,
input wire [44:0] MT_Layr_Minus_From_DataStream,
input wire MT_Layr_Minus_From_DataStream_en,
// Track Fits
output wire [125:0] CT_L1L2_DataStream,
output wire [125:0] CT_L3L4_DataStream,
output wire [125:0] CT_L5L6_DataStream,
output wire [125:0] CT_F1F2_DataStream,
output wire [125:0] CT_F3F4_DataStream,
output wire [125:0] CT_F1L1_DataStream

);

// Address bits "io_addr[31:30] = 2'b01" are consumed when selecting 'slave6'
// Address bits "io_addr[29:28] = 2'b01" are consumed when selecting 'tracklet_processing'
wire InputLink_R1Link1_io_sel, TPars_L1L2_io_sel;
wire InputLink_R1Link2_io_sel, TPars_L3L4_io_sel;
wire InputLink_R1Link3_io_sel, TPars_L5L6_io_sel;
wire io_sel_R3_io_block;
assign InputLink_R1Link1_io_sel = io_sel && (io_addr[13:10] == 4'b0001);
assign InputLink_R1Link2_io_sel = io_sel && (io_addr[13:10] == 4'b0010);
assign InputLink_R1Link3_io_sel = io_sel && (io_addr[13:10] == 4'b0011);
assign TPars_L1L2_io_sel  = io_sel && (io_addr[13:10] == 4'b0100);
assign TPars_L3L4_io_sel  = io_sel && (io_addr[13:10] == 4'b0101);
assign TPars_L5L6_io_sel  = io_sel && (io_addr[13:10] == 4'b0110);
assign io_sel_R3_io_block = io_sel && (io_addr[13:10] == 4'b1000);
// data busses for readback
wire [31:0] InputLink_R1Link1_io_rd_data, TPars_L1L2_io_rd_data;
wire [31:0] InputLink_R1Link2_io_rd_data, TPars_L3L4_io_rd_data;
wire [31:0] InputLink_R1Link3_io_rd_data, TPars_L5L6_io_rd_data;

wire IL1_D3_LR1_D3_empty;
wire IL2_D3_LR2_D3_empty;
wire IL3_D3_LR3_D3_empty;

reg [5:0] clk_cnt;

//wire enable_gen;
//enable_generator en_gen(
//.clk(clk),
//.in( (~IL1_D3_LR1_D3_empty | ~IL2_D3_LR2_D3_empty | ~IL3_D3_LR3_D3_empty) & bc0_i ),
//.out(enable_gen)
//);

initial
clk_cnt = 6'b0;
always @(posedge clk) begin
if(en_proc)
clk_cnt <= clk_cnt + 1'b1;
else begin
clk_cnt <= 6'b0;
end
if(clk_cnt == (`tmux - 1'b1))
clk_cnt <= 6'b0;
end

wire [1:0] IL1_D3_start;
wire [1:0] IL2_D3_start;
wire [1:0] IL3_D3_start;
wire [1:0] IL1_D4_start;
wire [1:0] IL2_D4_start;
wire [1:0] IL3_D4_start;
wire [1:0] IL1_D5_start;
wire [1:0] IL2_D5_start;
wire [1:0] IL3_D5_start;
wire [1:0] IL1_D6_start;
wire [1:0] IL2_D6_start;
wire [1:0] IL3_D6_start;

assign IL1_D3_start[1] = reset;    // use the top bit of start as reset
assign IL1_D3_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL2_D3_start[1] = reset;    // use the top bit of start as reset
assign IL2_D3_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL3_D3_start[1] = reset;    // use the top bit of start as reset
assign IL3_D3_start[0] = (clk_cnt == 6'd0 && en_proc);

assign IL1_D4_start[1] = reset;    // use the top bit of start as reset
assign IL1_D4_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL2_D4_start[1] = reset;    // use the top bit of start as reset
assign IL2_D4_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL3_D4_start[1] = reset;    // use the top bit of start as reset
assign IL3_D4_start[0] = (clk_cnt == 6'd0 && en_proc);

assign IL1_D5_start[1] = reset;    // use the top bit of start as reset
assign IL1_D5_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL2_D5_start[1] = reset;    // use the top bit of start as reset
assign IL2_D5_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL3_D5_start[1] = reset;    // use the top bit of start as reset
assign IL3_D5_start[0] = (clk_cnt == 6'd0 && en_proc);

assign IL1_D6_start[1] = reset;    // use the top bit of start as reset
assign IL1_D6_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL2_D6_start[1] = reset;    // use the top bit of start as reset
assign IL2_D6_start[0] = (clk_cnt == 6'd0 && en_proc);
assign IL3_D6_start[1] = reset;    // use the top bit of start as reset
assign IL3_D6_start[0] = (clk_cnt == 6'd0 && en_proc);


wire [1:0] TE_L3D3PHI2X2_L4D3PHI3X2_start;
wire [1:0] VMPROJ_L5L6_L1D3PHI2X2_start;
wire [1:0] PT_L3F3F5_Minus_start;
wire [1:0] VMPROJ_L1L2_L6D3PHI3X2_start;
wire [1:0] TPROJ_FromPlus_L4D4_L5L6_start;
wire [1:0] VMPROJ_L1L2_L3D4PHI3X1_start;
wire [1:0] VMPROJ_L5L6_L3D3PHI2X2_start;
wire [1:0] ME_L5L6_L4D3PHI2X2_start;
wire [1:0] TE_L5D4PHI3X2_L6D4PHI3X2_start;
wire [1:0] TE_L3D3PHI3X1_L4D3PHI3X2_start;
wire [1:0] PR_L4D4_L5L6_start;
wire [1:0] TE_L3D4PHI2X1_L4D4PHI2X1_start;
wire [1:0] VMPROJ_L3L4_L1D3PHI2X1_start;
wire [1:0] VMPROJ_L1L2_L5D4PHI3X2_start;
wire [1:0] ME_L5L6_L2D4PHI4X1_start;
wire [1:0] VMPROJ_L5L6_L4D3PHI2X2_start;
wire [1:0] VMS_L3D3PHI3X1n2_start;
wire [1:0] VMPROJ_L5L6_L3D4PHI2X2_start;
wire [1:0] ME_L3L4_L5D3PHI1X2_start;
wire [1:0] SP_L3D4PHI1X1_L4D4PHI1X1_start;
wire [1:0] ME_L3L4_L6D4PHI1X2_start;
wire [1:0] TE_L3D3PHI3X2_L4D3PHI3X2_start;
wire [1:0] VMS_L1D3PHI1X2n5_start;
wire [1:0] MC_L5L6_L1D4_start;
wire [1:0] ME_L3L4_L2D3PHI1X1_start;
wire [1:0] TE_L3D4PHI1X1_L4D4PHI1X2_start;
wire [1:0] ME_L5L6_L3D4PHI3X2_start;
wire [1:0] TE_L3D4PHI2X2_L4D4PHI2X2_start;
wire [1:0] VMPROJ_L1L2_L3D3PHI1X2_start;
wire [1:0] ME_L5L6_L1D4PHI2X1_start;
wire [1:0] SL1_L2D3_start;
wire [1:0] VMS_L1D3PHI3X1n6_start;
wire [1:0] VMPROJ_L5L6_L2D4PHI2X2_start;
wire [1:0] CM_L3L4_L1D3PHI1X1_start;
wire [1:0] VMS_L3D3PHI2X2n2_start;
wire [1:0] VMS_L5D4PHI2X1n3_start;
wire [1:0] VMPROJ_L5L6_L4D4PHI1X1_start;
wire [1:0] SP_L3D3PHI1X1_L4D3PHI1X1_start;
wire [1:0] VMS_L5D3PHI2X1n4_start;
wire [1:0] VMPROJ_L5L6_L4D3PHI3X2_start;
wire [1:0] TE_L1D4PHI3X1_L2D4PHI4X2_start;
wire [1:0] LR2_D4_start;
wire [1:0] VMR_L2D3_start;
wire [1:0] TE_L1D3PHI3X2_L2D4PHI4X2_start;
wire [1:0] VMPROJ_L3L4_L2D4PHI4X1_start;
wire [1:0] VMS_L1D3PHI3X1n4_start;
wire [1:0] VMS_L4D4PHI4X1n2_start;
wire [1:0] PR_L1D3_L3L4_start;
wire [1:0] TPROJ_FromPlus_L1D3_L3L4_start;
wire [1:0] TE_L1D3PHI1X1_L2D3PHI1X1_start;
wire [1:0] ME_L3L4_L6D3PHI1X1_start;
wire [1:0] ME_L5L6_L1D4PHI3X2_start;
wire [1:0] MC_L3L4_L1D4_start;
wire [1:0] PR_L2D3_L3L4_start;
wire [1:0] ME_L3L4_L2D4PHI3X2_start;
wire [1:0] CM_L3L4_L2D4PHI1X1_start;
wire [1:0] ME_L3L4_L6D3PHI2X2_start;
wire [1:0] VMS_L2D3PHI1X2n2_start;
wire [1:0] VMPROJ_L3L4_L5D4PHI3X2_start;
wire [1:0] TE_L3D4PHI1X2_L4D4PHI1X2_start;
wire [1:0] PR_L4D4_L1L2_start;
wire [1:0] MC_L3L4_L1D3_start;
wire [1:0] ME_L3L4_L6D3PHI3X2_start;
wire [1:0] MC_L3L4_L6D3_start;
wire [1:0] VMPROJ_L1L2_L5D4PHI2X2_start;
wire [1:0] VMPROJ_L3L4_L6D4PHI1X1_start;
wire [1:0] VMS_L2D4PHI2X2n3_start;
wire [1:0] VMPROJ_L3L4_L1D3PHI3X1_start;
wire [1:0] ME_L5L6_L2D4PHI1X1_start;
wire [1:0] ME_L1L2_L4D3PHI2X1_start;
wire [1:0] ME_L5L6_L4D4PHI4X2_start;
wire [1:0] ME_L1L2_L5D3PHI1X2_start;
wire [1:0] ME_L5L6_L4D4PHI2X2_start;
wire [1:0] TPROJ_ToMinus_L5D4L6D4_L1_start;
wire [1:0] FM_L5L6_L4_FromMinus_start;
wire [1:0] VMR_L6D4_start;
wire [1:0] VMPROJ_L3L4_L2D3PHI1X1_start;
wire [1:0] VMPROJ_L5L6_L4D3PHI4X2_start;
wire [1:0] VMS_L5D3PHI2X2n4_start;
wire [1:0] VMPROJ_L5L6_L4D4PHI4X1_start;
wire [1:0] VMPROJ_L1L2_L5D4PHI1X2_start;
wire [1:0] ME_L3L4_L5D3PHI1X1_start;
wire [1:0] VMS_L4D4PHI3X2n4_start;
wire [1:0] TE_L5D4PHI1X1_L6D4PHI2X2_start;
wire [1:0] ME_L1L2_L4D4PHI1X1_start;
wire [1:0] ME_L5L6_L3D3PHI1X2_start;
wire [1:0] SP_L1D4PHI1X1_L2D4PHI1X2_start;
wire [1:0] VMS_L1D3PHI3X1n5_start;
wire [1:0] VMPROJ_L1L2_L4D4PHI2X1_start;
wire [1:0] VMS_L3D3PHI1X2n1_start;
wire [1:0] LR3_D3_start;
wire [1:0] VMS_L5D4PHI2X1n4_start;
wire [1:0] ME_L5L6_L2D3PHI3X1_start;
wire [1:0] VMPROJ_L5L6_L1D3PHI2X1_start;
wire [1:0] TE_L1D3PHI3X2_L2D4PHI3X2_start;
wire [1:0] ME_L3L4_L6D4PHI3X1_start;
wire [1:0] VMPROJ_L5L6_L4D4PHI3X2_start;
wire [1:0] ME_L3L4_L2D3PHI4X1_start;
wire [1:0] VMR_L3D3_start;
wire [1:0] TE_L5D4PHI1X2_L6D4PHI2X2_start;
wire [1:0] TPROJ_FromPlus_L5D3_L3L4_start;
wire [1:0] VMPROJ_L1L2_L6D3PHI2X2_start;
wire [1:0] SL1_L3D4_start;
wire [1:0] VMS_L1D3PHI2X1n2_start;
wire [1:0] ME_L3L4_L2D4PHI4X2_start;
wire [1:0] VMS_L6D3PHI2X2n3_start;
wire [1:0] VMPROJ_L5L6_L4D4PHI2X2_start;
wire [1:0] TE_L5D4PHI3X1_L6D4PHI4X1_start;
wire [1:0] VMPROJ_L1L2_L4D3PHI2X1_start;
wire [1:0] CM_L5L6_L4D4PHI1X1_start;
wire [1:0] VMS_L3D4PHI2X1n4_start;
wire [1:0] SL1_L4D3_start;
wire [1:0] VMPROJ_L1L2_L5D3PHI1X2_start;
wire [1:0] SL1_L6D3_start;
wire [1:0] VMPROJ_L3L4_L2D3PHI1X2_start;
wire [1:0] ME_L3L4_L1D4PHI1X2_start;
wire [1:0] VMS_L6D3PHI1X2n2_start;
wire [1:0] ME_L1L2_L6D4PHI4X2_start;
wire [1:0] VMS_L2D4PHI2X2n4_start;
wire [1:0] TC_L5D4L6D4_proj_start;
wire [1:0] VMPROJ_L3L4_L2D3PHI4X2_start;
wire [1:0] TE_L3D3PHI2X2_L4D3PHI2X2_start;
wire [1:0] MC_L5L6_L4D4_start;
wire [1:0] TC_L1D4L2D4_start;
wire [1:0] PR_L4D3_L1L2_start;
wire [1:0] VMS_L4D4PHI3X1n3_start;
wire [1:0] TE_L5D3PHI2X2_L6D3PHI3X2_start;
wire [1:0] ME_L1L2_L3D4PHI2X1_start;
wire [1:0] ME_L1L2_L6D4PHI1X1_start;
wire [1:0] VMPROJ_L3L4_L1D3PHI1X2_start;
wire [1:0] PD_start;
wire [1:0] VMS_L5D4PHI3X1n4_start;
wire [1:0] VMPROJ_L5L6_L4D3PHI4X1_start;
wire [1:0] VMPROJ_L3L4_L2D3PHI4X1_start;
wire [1:0] MC_L1L2_L5D3_start;
wire [1:0] VMPROJ_L3L4_L6D3PHI3X2_start;
wire [1:0] TE_L5D4PHI2X2_L6D4PHI3X2_start;
wire [1:0] VMS_L1D3PHI1X2n4_start;
wire [1:0] SL1_L1D4_start;
wire [1:0] VMPROJ_L5L6_L4D4PHI3X1_start;
wire [1:0] TE_L1D3PHI3X1_L2D4PHI3X1_start;
wire [1:0] CM_L5L6_L3D4PHI1X1_start;
wire [1:0] VMPROJ_L1L2_L6D3PHI3X1_start;
wire [1:0] TE_L5D4PHI2X1_L6D4PHI2X2_start;
wire [1:0] VMPROJ_L5L6_L1D3PHI3X1_start;
wire [1:0] VMPROJ_L3L4_L1D3PHI3X2_start;
wire [1:0] MC_L1L2_L6D3_start;
wire [1:0] TC_L1D4L2D4_proj_start;
wire [1:0] ME_L5L6_L3D3PHI2X2_start;
wire [1:0] VMPROJ_L3L4_L1D4PHI2X1_start;
wire [1:0] ME_L5L6_L1D4PHI2X2_start;
wire [1:0] VMS_L5D3PHI2X1n3_start;
wire [1:0] ME_L3L4_L6D4PHI2X1_start;
wire [1:0] VMPROJ_L1L2_L6D3PHI1X1_start;
wire [1:0] VMPROJ_L5L6_L1D3PHI1X2_start;
wire [1:0] ME_L1L2_L5D3PHI3X1_start;
wire [1:0] PR_L6D3_L3L4_start;
wire [1:0] VMPROJ_L1L2_L4D4PHI3X1_start;
wire [1:0] VMS_L5D3PHI1X2n3_start;
wire [1:0] ME_L3L4_L6D4PHI4X2_start;
wire [1:0] VMPROJ_L5L6_L1D4PHI1X1_start;
wire [1:0] ME_L3L4_L5D4PHI3X2_start;
wire [1:0] VMPROJ_L5L6_L4D4PHI2X1_start;
wire [1:0] MC_L3L4_L5D3_start;
wire [1:0] VMS_L2D3PHI2X2n3_start;
wire [1:0] MC_L5L6_L3D3_start;
wire [1:0] VMPROJ_L3L4_L2D4PHI3X2_start;
wire [1:0] VMS_L5D3PHI3X1n4_start;
wire [1:0] VMS_L4D3PHI3X1n2_start;
wire [1:0] VMS_L1D3PHI3X2n5_start;
wire [1:0] VMPROJ_L5L6_L3D3PHI1X1_start;
wire [1:0] CM_L1L2_L3D4PHI1X1_start;
wire [1:0] VMPROJ_L3L4_L2D4PHI1X1_start;
wire [1:0] VMPROJ_L5L6_L4D3PHI3X1_start;
wire [1:0] VMS_L1D3PHI1X2n6_start;
wire [1:0] TE_L1D3PHI1X1_L2D3PHI2X2_start;
wire [1:0] TE_L5D3PHI3X2_L6D4PHI4X1_start;
wire [1:0] VMPROJ_L5L6_L3D3PHI1X2_start;
wire [1:0] VMS_L2D3PHI4X2n2_start;
wire [1:0] TPROJ_FromPlus_L3D4_L1L2_start;
wire [1:0] SP_L5D3PHI1X1_L6D3PHI1X1_start;
wire [1:0] SL1_L5D3_start;
wire [1:0] VMR_L3D4_start;
wire [1:0] TE_L1D3PHI3X2_L2D3PHI3X2_start;
wire [1:0] TE_L5D3PHI1X2_L6D4PHI2X1_start;
wire [1:0] TE_L3D3PHI3X1_L4D3PHI4X2_start;
wire [1:0] PR_L1D4_L5L6_start;
wire [1:0] TE_L5D4PHI1X1_L6D4PHI2X1_start;
wire [1:0] ME_L5L6_L1D4PHI3X1_start;
wire [1:0] VMPROJ_L1L2_L4D4PHI1X1_start;
wire [1:0] ME_L1L2_L6D4PHI4X1_start;
wire [1:0] FM_L3L4_L6_FromPlus_start;
wire [1:0] TE_L1D3PHI2X1_L2D3PHI2X2_start;
wire [1:0] TE_L1D3PHI2X1_L2D4PHI3X1_start;
wire [1:0] TC_L5D3L6D3_proj_start;
wire [1:0] TE_L5D3PHI1X1_L6D3PHI1X2_start;
wire [1:0] VMPROJ_L5L6_L2D4PHI4X2_start;
wire [1:0] VMPROJ_L3L4_L2D4PHI1X2_start;
wire [1:0] VMPROJ_L3L4_L1D4PHI3X2_start;
wire [1:0] TE_L1D3PHI1X1_L2D3PHI2X1_start;
wire [1:0] ME_L1L2_L6D3PHI1X2_start;
wire [1:0] VMPROJ_L1L2_L4D3PHI3X1_start;
wire [1:0] VMPROJ_L1L2_L6D4PHI3X2_start;
wire [1:0] VMPROJ_L5L6_L3D3PHI3X1_start;
wire [1:0] MC_L5L6_L2D4_start;
wire [1:0] VMS_L1D3PHI1X1n5_start;
wire [1:0] VMPROJ_L5L6_L2D3PHI3X1_start;
wire [1:0] VMPROJ_L3L4_L1D4PHI2X2_start;
wire [1:0] VMS_L3D3PHI1X1n4_start;
wire [1:0] ME_L1L2_L4D4PHI2X1_start;
wire [1:0] TE_L5D3PHI2X1_L6D3PHI3X1_start;
wire [1:0] TE_L3D3PHI2X1_L4D3PHI2X1_start;
wire [1:0] TE_L1D3PHI2X2_L2D4PHI2X1_start;
wire [1:0] SP_L3D3PHI1X2_L4D4PHI1X1_start;
wire [1:0] ME_L1L2_L5D3PHI3X2_start;
wire [1:0] CM_L1L2_L6D4PHI1X1_start;
wire [1:0] VMS_L3D4PHI1X1n4_start;
wire [1:0] ME_L5L6_L2D3PHI1X1_start;
wire [1:0] ME_L5L6_L4D4PHI1X1_start;
wire [1:0] VMS_L3D3PHI1X1n3_start;
wire [1:0] ME_L1L2_L5D4PHI1X2_start;
wire [1:0] ME_L3L4_L2D3PHI3X2_start;
wire [1:0] ME_L5L6_L3D4PHI2X2_start;
wire [1:0] TE_L1D3PHI2X2_L2D4PHI2X2_start;
wire [1:0] VMS_L1D3PHI1X1n6_start;
wire [1:0] VMS_L2D3PHI3X2n4_start;
wire [1:0] VMPROJ_L5L6_L4D4PHI1X2_start;
wire [1:0] ME_L5L6_L4D4PHI3X2_start;
wire [1:0] TE_L1D3PHI1X2_L2D4PHI2X1_start;
wire [1:0] VMPROJ_L5L6_L1D4PHI3X1_start;
wire [1:0] TE_L3D3PHI2X1_L4D3PHI3X2_start;
wire [1:0] VMS_L5D3PHI1X2n4_start;
wire [1:0] ME_L3L4_L1D4PHI3X2_start;
wire [1:0] ME_L5L6_L3D4PHI3X1_start;
wire [1:0] ME_L5L6_L2D4PHI2X2_start;
wire [1:0] TE_L1D4PHI2X1_L2D4PHI2X2_start;
wire [1:0] VMPROJ_L5L6_L1D4PHI2X1_start;
wire [1:0] VMS_L2D4PHI3X2n4_start;
wire [1:0] ME_L3L4_L5D4PHI2X2_start;
wire [1:0] LR1_D4_start;
wire [1:0] ME_L5L6_L2D3PHI2X1_start;
wire [1:0] VMR_L1D4_start;
wire [1:0] PR_L5D4_L1L2_start;
wire [1:0] TPROJ_ToPlus_L5D4L6D4_L1_start;
wire [1:0] TPROJ_FromPlus_L3D4_L5L6_start;
wire [1:0] VMPROJ_L5L6_L2D3PHI1X2_start;
wire [1:0] ME_L3L4_L5D4PHI3X1_start;
wire [1:0] TC_L5D3L6D4_proj_start;
wire [1:0] VMS_L3D3PHI1X2n3_start;
wire [1:0] ME_L5L6_L1D3PHI3X2_start;
wire [1:0] ME_L5L6_L3D4PHI1X2_start;
wire [1:0] ME_L5L6_L3D3PHI2X1_start;
wire [1:0] ME_L1L2_L5D4PHI2X2_start;
wire [1:0] MC_L5L6_L4D3_start;
wire [1:0] TE_L3D4PHI3X1_L4D4PHI4X2_start;
wire [1:0] TE_L1D3PHI2X2_L2D3PHI2X2_start;
wire [1:0] VMPROJ_L3L4_L5D3PHI3X1_start;
wire [1:0] TPROJ_ToPlus_L3D4L4D4_L5_start;
wire [1:0] TE_L5D3PHI1X2_L6D4PHI1X1_start;
wire [1:0] ME_L5L6_L2D4PHI3X2_start;
wire [1:0] PT_F1L5_Minus_start;
wire [1:0] VMS_L5D3PHI1X1n1_start;
wire [1:0] ME_L3L4_L6D4PHI1X1_start;
wire [1:0] VMS_L4D4PHI1X2n2_start;
wire [1:0] TPROJ_FromPlus_L6D4_L1L2_start;
wire [1:0] VMS_L1D3PHI2X2n6_start;
wire [1:0] TPROJ_ToMinus_L5D4L6D4_L4_start;
wire [1:0] ME_L1L2_L3D4PHI3X2_start;
wire [1:0] VMS_L6D3PHI4X2n2_start;
wire [1:0] ME_L1L2_L6D4PHI2X1_start;
wire [1:0] ME_L3L4_L6D4PHI4X1_start;
wire [1:0] MC_L3L4_L2D4_start;
wire [1:0] VMPROJ_L3L4_L6D4PHI4X1_start;
wire [1:0] CM_L3L4_L5D3PHI1X1_start;
wire [1:0] VMS_L2D3PHI3X2n3_start;
wire [1:0] VMPROJ_L3L4_L6D3PHI2X1_start;
wire [1:0] FT_L1L2_start;
wire [1:0] TE_L5D4PHI2X1_L6D4PHI3X2_start;
wire [1:0] ME_L3L4_L1D3PHI3X1_start;
wire [1:0] TE_L1D3PHI2X2_L2D4PHI3X1_start;
wire [1:0] ME_L3L4_L6D3PHI4X1_start;
wire [1:0] VMPROJ_L1L2_L3D3PHI2X1_start;
wire [1:0] CM_L3L4_L5D4PHI1X1_start;
wire [1:0] VMPROJ_L1L2_L3D3PHI3X2_start;
wire [1:0] ME_L5L6_L4D4PHI3X1_start;
wire [1:0] VMS_L1D3PHI3X1n3_start;
wire [1:0] ME_L1L2_L5D4PHI2X1_start;
wire [1:0] TE_L1D3PHI1X2_L2D4PHI2X2_start;
wire [1:0] MC_L1L2_L3D3_start;
wire [1:0] ME_L3L4_L1D3PHI1X2_start;
wire [1:0] TE_L5D3PHI1X1_L6D3PHI2X1_start;
wire [1:0] VMS_L3D3PHI3X2n2_start;
wire [1:0] VMS_L1D3PHI1X1n2_start;
wire [1:0] TE_L5D3PHI3X2_L6D4PHI3X1_start;
wire [1:0] ME_L5L6_L3D3PHI1X1_start;
wire [1:0] ME_L5L6_L4D3PHI2X1_start;
wire [1:0] VMS_L3D3PHI2X2n4_start;
wire [1:0] VMPROJ_L1L2_L5D3PHI3X2_start;
wire [1:0] VMPROJ_L1L2_L3D4PHI2X1_start;
wire [1:0] VMPROJ_L1L2_L5D3PHI2X2_start;
wire [1:0] VMS_L3D3PHI1X2n2_start;
wire [1:0] VMPROJ_L3L4_L6D3PHI2X2_start;
wire [1:0] TE_L3D3PHI3X2_L4D4PHI4X1_start;
wire [1:0] VMPROJ_L5L6_L3D4PHI3X2_start;
wire [1:0] VMPROJ_L1L2_L5D4PHI3X1_start;
wire [1:0] SP_L1D3PHI1X1_L2D4PHI1X1_start;
wire [1:0] TE_L3D4PHI2X1_L4D4PHI2X2_start;
wire [1:0] VMPROJ_L3L4_L5D4PHI1X2_start;
wire [1:0] VMS_L1D3PHI2X2n5_start;
wire [1:0] TE_L5D4PHI1X1_L6D4PHI1X1_start;
wire [1:0] VMPROJ_L1L2_L5D4PHI2X1_start;
wire [1:0] VMPROJ_L3L4_L2D4PHI4X2_start;
wire [1:0] TE_L3D3PHI2X2_L4D4PHI3X1_start;
wire [1:0] ME_L5L6_L1D4PHI1X1_start;
wire [1:0] ME_L3L4_L1D4PHI2X1_start;
wire [1:0] TC_L1D3L2D4_start;
wire [1:0] ME_L5L6_L3D3PHI3X1_start;
wire [1:0] VMS_L1D3PHI2X2n3_start;
wire [1:0] VMPROJ_L1L2_L3D4PHI2X2_start;
wire [1:0] TE_L3D4PHI3X2_L4D4PHI4X2_start;
wire [1:0] VMPROJ_L5L6_L1D4PHI2X2_start;
wire [1:0] TE_L3D4PHI3X2_L4D4PHI3X2_start;
wire [1:0] TE_L3D4PHI1X1_L4D4PHI2X2_start;
wire [1:0] CM_L3L4_L6D3PHI1X1_start;
wire [1:0] TE_L1D3PHI2X1_L2D4PHI2X1_start;
wire [1:0] ME_L1L2_L3D3PHI3X1_start;
wire [1:0] VMPROJ_L1L2_L5D4PHI1X1_start;
wire [1:0] VMS_L5D3PHI2X2n3_start;
wire [1:0] VMPROJ_L5L6_L3D4PHI2X1_start;
wire [1:0] VMPROJ_L5L6_L2D4PHI3X2_start;
wire [1:0] VMPROJ_L5L6_L3D3PHI2X1_start;
wire [1:0] VMS_L6D4PHI3X1n4_start;
wire [1:0] ME_L1L2_L4D4PHI1X2_start;
wire [1:0] PR_L6D4_L1L2_start;
wire [1:0] VMPROJ_L5L6_L3D4PHI1X1_start;
wire [1:0] ME_L1L2_L6D3PHI1X1_start;
wire [1:0] TPROJ_FromPlus_L5D4_L3L4_start;
wire [1:0] ME_L5L6_L4D3PHI1X2_start;
wire [1:0] TE_L3D3PHI2X1_L4D3PHI2X2_start;
wire [1:0] VMPROJ_L3L4_L1D4PHI1X1_start;
wire [1:0] ME_L3L4_L2D4PHI3X1_start;
wire [1:0] ME_L3L4_L6D4PHI3X2_start;
wire [1:0] MC_L1L2_L6D4_start;
wire [1:0] VMS_L1D3PHI2X1n5_start;
wire [1:0] VMS_L5D3PHI3X2n4_start;
wire [1:0] ME_L1L2_L4D3PHI4X2_start;
wire [1:0] VMS_L3D4PHI1X1n3_start;
wire [1:0] ME_L5L6_L2D3PHI4X2_start;
wire [1:0] PR_L4D3_L5L6_start;
wire [1:0] VMS_L3D3PHI3X1n3_start;
wire [1:0] VMS_L4D4PHI4X2n2_start;
wire [1:0] VMS_L4D4PHI2X1n4_start;
wire [1:0] VMS_L6D4PHI3X2n3_start;
wire [1:0] TE_L3D3PHI1X2_L4D3PHI2X2_start;
wire [1:0] VMPROJ_L3L4_L6D4PHI1X2_start;
wire [1:0] ME_L1L2_L3D3PHI2X2_start;
wire [1:0] VMPROJ_L3L4_L5D4PHI3X1_start;
wire [1:0] VMPROJ_L1L2_L6D4PHI1X1_start;
wire [1:0] PT_L1L6F4_Minus_start;
wire [1:0] TE_L5D3PHI2X2_L6D4PHI2X1_start;
wire [1:0] ME_L1L2_L5D3PHI2X1_start;
wire [1:0] ME_L5L6_L1D3PHI3X1_start;
wire [1:0] VMPROJ_L3L4_L1D4PHI3X1_start;
wire [1:0] VMS_L3D3PHI3X2n4_start;
wire [1:0] TE_L5D4PHI3X1_L6D4PHI4X2_start;
wire [1:0] ME_L5L6_L1D4PHI1X2_start;
wire [1:0] MC_L5L6_L2D3_start;
wire [1:0] VMS_L2D4PHI4X2n2_start;
wire [1:0] TPROJ_ToPlus_L5D4L6D4_L4_start;
wire [1:0] ME_L1L2_L4D3PHI1X1_start;
wire [1:0] VMS_L1D3PHI3X2n6_start;
wire [1:0] TE_L5D3PHI1X2_L6D3PHI2X2_start;
wire [1:0] ME_L1L2_L5D4PHI3X1_start;
wire [1:0] CM_L1L2_L4D4PHI1X1_start;
wire [1:0] ME_L5L6_L2D4PHI4X2_start;
wire [1:0] PT_F1L5_Plus_start;
wire [1:0] PR_L3D3_L1L2_start;
wire [1:0] ME_L3L4_L5D4PHI1X2_start;
wire [1:0] VMS_L1D3PHI3X2n3_start;
wire [1:0] SP_L1D3PHI1X1_L2D3PHI1X1_start;
wire [1:0] ME_L1L2_L5D3PHI2X2_start;
wire [1:0] ME_L5L6_L4D4PHI4X1_start;
wire [1:0] TC_L1D3L2D4_proj_start;
wire [1:0] FM_L1L2_L3D3_ToPlus_start;
wire [1:0] TE_L3D3PHI2X1_L4D3PHI3X1_start;
wire [1:0] ME_L1L2_L6D3PHI4X1_start;
wire [1:0] VMS_L5D3PHI3X1n2_start;
wire [1:0] MT_Layr_Plus_start;
wire [1:0] SL1_L1D3_start;
wire [1:0] TE_L1D3PHI1X1_L2D4PHI2X1_start;
wire [1:0] MC_L3L4_L6D4_start;
wire [1:0] ME_L1L2_L6D4PHI3X1_start;
wire [1:0] ME_L5L6_L4D4PHI2X1_start;
wire [1:0] VMPROJ_L3L4_L1D3PHI2X2_start;
wire [1:0] TE_L5D4PHI3X1_L6D4PHI3X2_start;
wire [1:0] ME_L5L6_L2D3PHI3X2_start;
wire [1:0] TE_L1D3PHI2X1_L2D3PHI3X1_start;
wire [1:0] ME_L3L4_L1D3PHI2X1_start;
wire [1:0] ME_L3L4_L5D3PHI3X1_start;
wire [1:0] ME_L5L6_L2D3PHI1X2_start;
wire [1:0] TE_L5D3PHI2X2_L6D3PHI2X2_start;
wire [1:0] ME_L3L4_L2D3PHI4X2_start;
wire [1:0] VMS_L5D3PHI3X2n3_start;
wire [1:0] ME_L3L4_L2D4PHI4X1_start;
wire [1:0] ME_L5L6_L1D3PHI1X1_start;
wire [1:0] VMS_L4D3PHI2X1n2_start;
wire [1:0] PR_L5D3_L3L4_start;
wire [1:0] ME_L1L2_L4D3PHI3X1_start;
wire [1:0] SL1_L2D4_start;
wire [1:0] TPROJ_FromPlus_L2D3_L5L6_start;
wire [1:0] ME_L1L2_L5D4PHI3X2_start;
wire [1:0] VMPROJ_L3L4_L5D3PHI2X1_start;
wire [1:0] ME_L3L4_L6D3PHI3X1_start;
wire [1:0] TC_L5D3L6D3_start;
wire [1:0] FT_L5L6_start;
wire [1:0] LR1_D3_start;
wire [1:0] VMS_L3D3PHI1X1n1_start;
wire [1:0] TPROJ_FromPlus_L4D3_L5L6_start;
wire [1:0] VMPROJ_L3L4_L6D3PHI1X2_start;
wire [1:0] VMS_L1D3PHI3X2n4_start;
wire [1:0] VMPROJ_L3L4_L1D4PHI1X2_start;
wire [1:0] ME_L3L4_L2D3PHI3X1_start;
wire [1:0] TPROJ_FromPlus_L2D3_L3L4_start;
wire [1:0] ME_L1L2_L3D4PHI1X1_start;
wire [1:0] VMR_L4D4_start;
wire [1:0] MC_L1L2_L3D4_start;
wire [1:0] ME_L3L4_L2D3PHI2X2_start;
wire [1:0] TE_L5D3PHI2X2_L6D4PHI3X1_start;
wire [1:0] VMS_L4D4PHI2X1n3_start;
wire [1:0] VMPROJ_L3L4_L2D3PHI2X2_start;
wire [1:0] VMPROJ_L1L2_L4D3PHI1X2_start;
wire [1:0] TPROJ_FromPlus_L2D4_L3L4_start;
wire [1:0] TC_L1D3L2D3_proj_start;
wire [1:0] ME_L3L4_L1D3PHI3X2_start;
wire [1:0] VMPROJ_L3L4_L1D3PHI1X1_start;
wire [1:0] VMPROJ_L3L4_L2D3PHI3X1_start;
wire [1:0] VMS_L6D3PHI3X1n2_start;
wire [1:0] VMPROJ_L3L4_L6D4PHI3X1_start;
wire [1:0] VMS_L6D4PHI2X1n3_start;
wire [1:0] ME_L1L2_L6D4PHI1X2_start;
wire [1:0] VMPROJ_L1L2_L3D4PHI1X2_start;
wire [1:0] VMPROJ_L5L6_L1D4PHI3X2_start;
wire [1:0] ME_L3L4_L2D4PHI1X1_start;
wire [1:0] TE_L1D3PHI1X1_L2D3PHI1X2_start;
wire [1:0] VMPROJ_L1L2_L6D3PHI1X2_start;
wire [1:0] VMS_L5D3PHI1X1n2_start;
wire [1:0] VMS_L5D3PHI2X1n2_start;
wire [1:0] TE_L5D4PHI2X1_L6D4PHI2X1_start;
wire [1:0] ME_L1L2_L4D4PHI4X1_start;
wire [1:0] TPROJ_FromPlus_L6D3_L3L4_start;
wire [1:0] ME_L1L2_L4D4PHI3X1_start;
wire [1:0] VMS_L1D3PHI2X1n4_start;
wire [1:0] ME_L5L6_L2D3PHI4X1_start;
wire [1:0] ME_L1L2_L6D3PHI3X2_start;
wire [1:0] MC_L3L4_L5D4_start;
wire [1:0] VMPROJ_L1L2_L4D4PHI3X2_start;
wire [1:0] VMPROJ_L1L2_L6D3PHI4X1_start;
wire [1:0] VMPROJ_L1L2_L6D4PHI1X2_start;
wire [1:0] ME_L5L6_L1D3PHI2X2_start;
wire [1:0] TC_L3D3L4D4_start;
wire [1:0] VMPROJ_L1L2_L6D4PHI4X2_start;
wire [1:0] VMPROJ_L5L6_L2D4PHI4X1_start;
wire [1:0] ME_L1L2_L3D4PHI1X2_start;
wire [1:0] VMPROJ_L5L6_L1D4PHI1X2_start;
wire [1:0] VMPROJ_L5L6_L2D3PHI1X1_start;
wire [1:0] ME_L3L4_L6D3PHI4X2_start;
wire [1:0] VMS_L6D3PHI3X2n4_start;
wire [1:0] VMPROJ_L1L2_L6D4PHI4X1_start;
wire [1:0] VMPROJ_L3L4_L5D3PHI1X2_start;
wire [1:0] ME_L3L4_L1D4PHI1X1_start;
wire [1:0] VMS_L4D4PHI2X2n3_start;
wire [1:0] TE_L5D4PHI3X1_L6D4PHI3X1_start;
wire [1:0] TE_L1D3PHI3X1_L2D3PHI4X2_start;
wire [1:0] VMPROJ_L3L4_L5D3PHI1X1_start;
wire [1:0] CM_L5L6_L1D3PHI1X1_start;
wire [1:0] TE_L3D3PHI3X1_L4D3PHI4X1_start;
wire [1:0] MC_L1L2_L4D3_start;
wire [1:0] TE_L3D4PHI3X1_L4D4PHI4X1_start;
wire [1:0] ME_L1L2_L6D3PHI2X1_start;
wire [1:0] TE_L3D4PHI1X2_L4D4PHI2X2_start;
wire [1:0] TC_L1D3L2D3_start;
wire [1:0] PR_L2D4_L5L6_start;
wire [1:0] VMS_L1D3PHI2X1n6_start;
wire [1:0] TE_L1D3PHI2X2_L2D3PHI3X2_start;
wire [1:0] TE_L3D3PHI1X1_L4D3PHI2X1_start;
wire [1:0] VMR_L2D4_start;
wire [1:0] PR_L1D3_L5L6_start;
wire [1:0] VMS_L4D3PHI3X2n2_start;
wire [1:0] VMPROJ_L1L2_L5D3PHI3X1_start;
wire [1:0] VMPROJ_L5L6_L1D3PHI1X1_start;
wire [1:0] TE_L3D4PHI3X1_L4D4PHI3X1_start;
wire [1:0] TPROJ_FromPlus_L1D4_L3L4_start;
wire [1:0] SL1_L4D4_start;
wire [1:0] VMPROJ_L1L2_L3D3PHI1X1_start;
wire [1:0] ME_L3L4_L5D3PHI2X1_start;
wire [1:0] TE_L5D3PHI1X1_L6D3PHI2X2_start;
wire [1:0] TPROJ_FromPlus_L1D3_L5L6_start;
wire [1:0] ME_L3L4_L2D3PHI1X2_start;
wire [1:0] TE_L1D4PHI1X1_L2D4PHI2X2_start;
wire [1:0] VMPROJ_L5L6_L1D3PHI3X2_start;
wire [1:0] TE_L3D4PHI1X1_L4D4PHI1X1_start;
wire [1:0] ME_L1L2_L4D3PHI1X2_start;
wire [1:0] VMS_L1D3PHI1X1n1_start;
wire [1:0] ME_L3L4_L2D4PHI1X2_start;
wire [1:0] CM_L3L4_L6D4PHI1X1_start;
wire [1:0] VMS_L6D4PHI1X2n2_start;
wire [1:0] ME_L1L2_L6D3PHI3X1_start;
wire [1:0] MC_L5L6_L1D3_start;
wire [1:0] PR_L5D4_L3L4_start;
wire [1:0] TE_L3D3PHI3X2_L4D3PHI4X2_start;
wire [1:0] VMPROJ_L1L2_L4D4PHI4X1_start;
wire [1:0] TE_L3D3PHI3X2_L4D4PHI3X1_start;
wire [1:0] ME_L1L2_L3D3PHI2X1_start;
wire [1:0] VMS_L1D3PHI2X2n4_start;
wire [1:0] TE_L1D3PHI3X1_L2D3PHI3X1_start;
wire [1:0] TE_L1D3PHI1X2_L2D4PHI1X2_start;
wire [1:0] TE_L5D3PHI3X1_L6D3PHI4X2_start;
wire [1:0] PR_L5D3_L1L2_start;
wire [1:0] TPROJ_ToMinus_L5D4L6D4_L3_start;
wire [1:0] ME_L1L2_L4D4PHI4X2_start;
wire [1:0] VMS_L4D3PHI2X2n2_start;
wire [1:0] ME_L1L2_L5D3PHI1X1_start;
wire [1:0] VMPROJ_L5L6_L2D3PHI4X2_start;
wire [1:0] VMS_L5D4PHI1X1n3_start;
wire [1:0] CM_L5L6_L2D3PHI1X1_start;
wire [1:0] VMS_L3D3PHI3X1n4_start;
wire [1:0] TPROJ_ToPlus_L5D4L6D4_L3_start;
wire [1:0] VMS_L1D3PHI1X2n3_start;
wire [1:0] ME_L5L6_L2D4PHI1X2_start;
wire [1:0] VMS_L5D4PHI3X1n3_start;
wire [1:0] VMS_L4D4PHI1X1n2_start;
wire [1:0] VMS_L1D3PHI3X1n2_start;
wire [1:0] ME_L3L4_L5D3PHI2X2_start;
wire [1:0] TE_L3D3PHI2X2_L4D4PHI2X1_start;
wire [1:0] TE_L3D4PHI2X1_L4D4PHI3X2_start;
wire [1:0] VMPROJ_L1L2_L4D3PHI4X1_start;
wire [1:0] ME_L1L2_L5D4PHI1X1_start;
wire [1:0] VMS_L6D4PHI1X1n2_start;
wire [1:0] TE_L3D3PHI1X2_L4D4PHI2X1_start;
wire [1:0] VMPROJ_L1L2_L4D3PHI2X2_start;
wire [1:0] SL1_L6D4_start;
wire [1:0] TE_L1D3PHI2X2_L2D4PHI3X2_start;
wire [1:0] LR3_D4_start;
wire [1:0] TC_L5D3L6D4_start;
wire [1:0] TE_L5D3PHI3X1_L6D3PHI3X1_start;
wire [1:0] VMPROJ_L3L4_L6D4PHI3X2_start;
wire [1:0] FM_L1L2_L3D3_ToMinus_start;
wire [1:0] TPROJ_ToMinus_L3D4L4D4_L5_start;
wire [1:0] ME_L5L6_L3D3PHI3X2_start;
wire [1:0] VMPROJ_L3L4_L6D3PHI3X1_start;
wire [1:0] VMS_L3D3PHI1X2n4_start;
wire [1:0] ME_L3L4_L5D4PHI2X1_start;
wire [1:0] TE_L5D4PHI1X2_L6D4PHI1X2_start;
wire [1:0] VMPROJ_L5L6_L3D3PHI3X2_start;
wire [1:0] PT_L1L6F4_Plus_start;
wire [1:0] TPROJ_FromPlus_L2D4_L5L6_start;
wire [1:0] TE_L1D3PHI3X1_L2D3PHI4X1_start;
wire [1:0] VMR_L5D3_start;
wire [1:0] MC_L1L2_L4D4_start;
wire [1:0] VMPROJ_L1L2_L6D4PHI3X1_start;
wire [1:0] VMS_L2D4PHI1X2n2_start;
wire [1:0] TE_L1D3PHI1X2_L2D4PHI1X1_start;
wire [1:0] VMPROJ_L3L4_L5D3PHI3X2_start;
wire [1:0] VMPROJ_L1L2_L5D3PHI1X1_start;
wire [1:0] ME_L3L4_L6D4PHI2X2_start;
wire [1:0] VMS_L3D3PHI2X1n2_start;
wire [1:0] PR_L2D3_L5L6_start;
wire [1:0] CM_L1L2_L6D3PHI1X1_start;
wire [1:0] TE_L3D3PHI1X1_L4D3PHI1X1_start;
wire [1:0] PR_L6D4_L3L4_start;
wire [1:0] VMS_L3D3PHI2X1n4_start;
wire [1:0] ME_L1L2_L6D3PHI2X2_start;
wire [1:0] TE_L5D3PHI1X1_L6D3PHI1X1_start;
wire [1:0] CM_L1L2_L3D3PHI1X1_start;
wire [1:0] VMPROJ_L3L4_L6D3PHI1X1_start;
wire [1:0] MT_Layr_Minus_start;
wire [1:0] VMS_L3D3PHI1X1n2_start;
wire [1:0] VMS_L5D3PHI1X1n4_start;
wire [1:0] VMPROJ_L1L2_L3D3PHI2X2_start;
wire [1:0] ME_L5L6_L2D4PHI2X1_start;
wire [1:0] ME_L1L2_L4D4PHI3X2_start;
wire [1:0] VMPROJ_L5L6_L2D4PHI1X2_start;
wire [1:0] MC_L1L2_L5D4_start;
wire [1:0] CM_L1L2_L4D3PHI1X1_start;
wire [1:0] ME_L1L2_L3D4PHI3X1_start;
wire [1:0] TPROJ_FromPlus_L5D4_L1L2_start;
wire [1:0] PR_L1D4_L3L4_start;
wire [1:0] TE_L3D4PHI3X1_L4D4PHI3X2_start;
wire [1:0] VMS_L3D3PHI2X2n3_start;
wire [1:0] VMPROJ_L5L6_L2D4PHI3X1_start;
wire [1:0] ME_L5L6_L4D3PHI3X1_start;
wire [1:0] VMPROJ_L3L4_L6D4PHI4X2_start;
wire [1:0] ME_L5L6_L4D3PHI4X1_start;
wire [1:0] VMPROJ_L5L6_L4D3PHI1X1_start;
wire [1:0] VMPROJ_L3L4_L5D4PHI2X1_start;
wire [1:0] TC_L3D4L4D4_proj_start;
wire [1:0] VMPROJ_L3L4_L2D4PHI3X1_start;
wire [1:0] VMS_L6D3PHI3X2n3_start;
wire [1:0] VMS_L4D4PHI3X2n3_start;
wire [1:0] ME_L3L4_L6D3PHI1X2_start;
wire [1:0] VMS_L5D3PHI1X1n3_start;
wire [1:0] PR_L3D3_L5L6_start;
wire [1:0] TC_L5D4L6D4_start;
wire [1:0] PR_L3D4_L5L6_start;
wire [1:0] ME_L1L2_L3D3PHI1X1_start;
wire [1:0] ME_L5L6_L4D3PHI1X1_start;
wire [1:0] VMS_L1D3PHI1X1n3_start;
wire [1:0] VMPROJ_L1L2_L3D3PHI3X1_start;
wire [1:0] VMS_L2D3PHI2X1n2_start;
wire [1:0] ME_L1L2_L4D3PHI4X1_start;
wire [1:0] VMS_L6D3PHI2X1n2_start;
wire [1:0] ME_L5L6_L3D4PHI1X1_start;
wire [1:0] VMS_L6D4PHI3X2n4_start;
wire [1:0] VMPROJ_L5L6_L2D3PHI2X1_start;
wire [1:0] VMPROJ_L1L2_L3D4PHI3X2_start;
wire [1:0] TE_L1D3PHI3X2_L2D4PHI4X1_start;
wire [1:0] VMR_L4D3_start;
wire [1:0] VMPROJ_L5L6_L2D4PHI1X1_start;
wire [1:0] VMPROJ_L1L2_L4D4PHI2X2_start;
wire [1:0] TPROJ_FromPlus_L3D3_L1L2_start;
wire [1:0] TE_L3D3PHI3X1_L4D3PHI3X1_start;
wire [1:0] VMPROJ_L3L4_L6D4PHI2X1_start;
wire [1:0] ME_L1L2_L3D4PHI2X2_start;
wire [1:0] CM_L5L6_L3D3PHI1X1_start;
wire [1:0] TE_L1D3PHI2X1_L2D3PHI2X1_start;
wire [1:0] CM_L5L6_L4D3PHI1X1_start;
wire [1:0] TE_L5D4PHI1X1_L6D4PHI1X2_start;
wire [1:0] TE_L1D3PHI3X1_L2D4PHI4X1_start;
wire [1:0] VMS_L6D4PHI4X1n2_start;
wire [1:0] TC_L3D4L4D4_start;
wire [1:0] VMPROJ_L3L4_L5D4PHI1X1_start;
wire [1:0] VMPROJ_L5L6_L2D3PHI3X2_start;
wire [1:0] VMPROJ_L1L2_L6D4PHI2X2_start;
wire [1:0] TC_L3D3L4D4_proj_start;
wire [1:0] ME_L3L4_L1D4PHI2X2_start;
wire [1:0] ME_L3L4_L1D4PHI3X1_start;
wire [1:0] TE_L1D3PHI1X1_L2D4PHI1X1_start;
wire [1:0] PR_L6D3_L1L2_start;
wire [1:0] VMS_L6D4PHI2X1n4_start;
wire [1:0] ME_L3L4_L2D4PHI2X1_start;
wire [1:0] SL1_L5D4_start;
wire [1:0] VMPROJ_L1L2_L4D4PHI1X2_start;
wire [1:0] TE_L1D3PHI3X2_L2D3PHI4X2_start;
wire [1:0] SL1_L3D3_start;
wire [1:0] TE_L1D4PHI3X1_L2D4PHI3X2_start;
wire [1:0] VMPROJ_L5L6_L4D3PHI2X1_start;
wire [1:0] TE_L3D4PHI2X2_L4D4PHI3X2_start;
wire [1:0] CM_L5L6_L1D4PHI1X1_start;
wire [1:0] TPROJ_FromPlus_L5D3_L1L2_start;
wire [1:0] PT_L2L4F2_Plus_start;
wire [1:0] TC_L3D3L4D3_proj_start;
wire [1:0] ME_L1L2_L6D4PHI3X2_start;
wire [1:0] ME_L1L2_L6D3PHI4X2_start;
wire [1:0] VMPROJ_L1L2_L6D4PHI2X1_start;
wire [1:0] TE_L5D4PHI2X2_L6D4PHI2X2_start;
wire [1:0] PT_L2L4F2_Minus_start;
wire [1:0] VMPROJ_L5L6_L2D4PHI2X1_start;
wire [1:0] VMPROJ_L3L4_L5D3PHI2X2_start;
wire [1:0] ME_L3L4_L1D3PHI2X2_start;
wire [1:0] TE_L3D4PHI1X1_L4D4PHI2X1_start;
wire [1:0] TE_L3D3PHI1X1_L4D3PHI1X2_start;
wire [1:0] TE_L1D3PHI1X2_L2D3PHI2X2_start;
wire [1:0] TE_L1D4PHI2X1_L2D4PHI3X2_start;
wire [1:0] TPROJ_FromPlus_L6D4_L3L4_start;
wire [1:0] ME_L1L2_L3D3PHI3X2_start;
wire [1:0] VMPROJ_L5L6_L2D3PHI4X1_start;
wire [1:0] VMS_L3D3PHI2X1n3_start;
wire [1:0] VMS_L3D4PHI3X1n4_start;
wire [1:0] ME_L5L6_L4D4PHI1X2_start;
wire [1:0] ME_L5L6_L4D3PHI3X2_start;
wire [1:0] VMPROJ_L5L6_L4D4PHI4X2_start;
wire [1:0] VMPROJ_L5L6_L2D3PHI2X2_start;
wire [1:0] VMPROJ_L3L4_L6D4PHI2X2_start;
wire [1:0] VMS_L2D3PHI3X1n2_start;
wire [1:0] TE_L3D3PHI1X2_L4D3PHI1X2_start;
wire [1:0] VMS_L6D4PHI2X2n3_start;
wire [1:0] SP_L5D4PHI1X1_L6D4PHI1X1_start;
wire [1:0] TPROJ_FromPlus_L6D3_L1L2_start;
wire [1:0] LR2_D3_start;
wire [1:0] TE_L5D3PHI3X2_L6D3PHI4X2_start;
wire [1:0] VMPROJ_L3L4_L2D3PHI3X2_start;
wire [1:0] ME_L1L2_L4D3PHI3X2_start;
wire [1:0] VMPROJ_L1L2_L3D4PHI1X1_start;
wire [1:0] VMPROJ_L1L2_L6D3PHI2X1_start;
wire [1:0] VMS_L3D3PHI3X2n3_start;
wire [1:0] TE_L3D3PHI1X2_L4D4PHI1X1_start;
wire [1:0] ME_L1L2_L3D3PHI1X2_start;
wire [1:0] TE_L5D3PHI2X1_L6D3PHI3X2_start;
wire [1:0] TPROJ_FromPlus_L4D3_L1L2_start;
wire [1:0] ME_L3L4_L2D3PHI2X1_start;
wire [1:0] VMR_L1D3_start;
wire [1:0] VMS_L1D3PHI2X1n3_start;
wire [1:0] TC_L3D3L4D3_start;
wire [1:0] CM_L3L4_L2D3PHI1X1_start;
wire [1:0] VMPROJ_L1L2_L4D3PHI4X2_start;
wire [1:0] ME_L1L2_L4D4PHI2X2_start;
wire [1:0] VMR_L5D4_start;
wire [1:0] VMPROJ_L1L2_L4D4PHI4X2_start;
wire [1:0] VMPROJ_L3L4_L2D4PHI2X1_start;
wire [1:0] TPROJ_FromPlus_L3D3_L5L6_start;
wire [1:0] ME_L5L6_L3D4PHI2X1_start;
wire [1:0] MC_L5L6_L3D4_start;
wire [1:0] ME_L1L2_L6D4PHI2X2_start;
wire [1:0] CM_L5L6_L2D4PHI1X1_start;
wire [1:0] ME_L5L6_L1D3PHI2X1_start;
wire [1:0] VMPROJ_L5L6_L4D3PHI1X2_start;
wire [1:0] TPROJ_FromPlus_L4D4_L1L2_start;
wire [1:0] VMPROJ_L5L6_L3D4PHI1X2_start;
wire [1:0] ME_L3L4_L5D4PHI1X1_start;
wire [1:0] SP_L5D3PHI1X2_L6D4PHI1X1_start;
wire [1:0] TE_L3D3PHI1X1_L4D3PHI2X2_start;
wire [1:0] VMS_L5D3PHI3X1n3_start;
wire [1:0] VMS_L6D4PHI3X1n3_start;
wire [1:0] ME_L3L4_L2D4PHI2X2_start;
wire [1:0] VMS_L2D4PHI3X2n3_start;
wire [1:0] TE_L1D3PHI3X1_L2D3PHI3X2_start;
wire [1:0] VMPROJ_L1L2_L4D3PHI1X1_start;
wire [1:0] ME_L3L4_L6D3PHI2X1_start;
wire [1:0] TPROJ_FromPlus_L1D4_L5L6_start;
wire [1:0] TE_L5D3PHI2X1_L6D3PHI2X1_start;
wire [1:0] VMR_L6D3_start;
wire [1:0] VMS_L5D4PHI1X1n4_start;
wire [1:0] TE_L1D3PHI1X2_L2D3PHI1X2_start;
wire [1:0] TE_L1D3PHI2X1_L2D3PHI3X2_start;
wire [1:0] TE_L3D4PHI2X1_L4D4PHI3X1_start;
wire [1:0] MC_L3L4_L2D3_start;
wire [1:0] TE_L1D4PHI1X1_L2D4PHI1X2_start;
wire [1:0] VMPROJ_L3L4_L2D4PHI2X2_start;
wire [1:0] ME_L5L6_L4D3PHI4X2_start;
wire [1:0] VMPROJ_L3L4_L5D4PHI2X2_start;
wire [1:0] CM_L1L2_L5D3PHI1X1_start;
wire [1:0] ME_L3L4_L1D3PHI1X1_start;
wire [1:0] TE_L5D3PHI1X2_L6D3PHI1X2_start;
wire [1:0] TE_L5D3PHI3X1_L6D3PHI4X1_start;
wire [1:0] TE_L5D4PHI3X2_L6D4PHI4X2_start;
wire [1:0] VMS_L4D4PHI3X1n4_start;
wire [1:0] TE_L5D3PHI3X1_L6D3PHI3X2_start;
wire [1:0] TE_L5D4PHI2X1_L6D4PHI3X1_start;
wire [1:0] CM_L1L2_L5D4PHI1X1_start;
wire [1:0] VMS_L3D4PHI2X1n3_start;
wire [1:0] VMS_L6D4PHI2X2n4_start;
wire [1:0] ME_L5L6_L2D4PHI3X1_start;
wire [1:0] ME_L1L2_L4D3PHI2X2_start;
wire [1:0] TE_L5D3PHI3X2_L6D3PHI3X2_start;
wire [1:0] TE_L1D3PHI3X2_L2D4PHI3X1_start;
wire [1:0] TE_L5D3PHI2X1_L6D3PHI2X2_start;
wire [1:0] FM_L1L2_L6_FromMinus_start;
wire [1:0] TF_L1L2_start;
wire [1:0] VMS_L6D3PHI2X2n4_start;
wire [1:0] VMPROJ_L5L6_L3D4PHI3X1_start;
wire [1:0] PT_L3F3F5_Plus_start;
wire [1:0] VMS_L6D4PHI4X2n2_start;
wire [1:0] FT_L3L4_start;
wire [1:0] CM_L3L4_L1D4PHI1X1_start;
wire [1:0] VMPROJ_L3L4_L6D3PHI4X1_start;
wire [1:0] VMPROJ_L3L4_L2D3PHI2X1_start;
wire [1:0] ME_L5L6_L2D3PHI2X2_start;
wire [1:0] VMS_L4D4PHI2X2n4_start;
wire [1:0] VMPROJ_L1L2_L5D3PHI2X1_start;
wire [1:0] ME_L3L4_L5D3PHI3X2_start;
wire [1:0] PR_L2D4_L3L4_start;
wire [1:0] VMS_L3D4PHI3X1n3_start;
wire [1:0] VMPROJ_L1L2_L4D3PHI3X2_start;
wire [1:0] VMPROJ_L3L4_L6D3PHI4X2_start;
wire [1:0] VMS_L2D3PHI2X2n4_start;
wire [1:0] VMPROJ_L1L2_L6D3PHI4X2_start;
wire [1:0] PR_L3D4_L1L2_start;
wire [1:0] ME_L5L6_L1D3PHI1X2_start;
wire [1:0] VMS_L1D3PHI1X1n4_start;

wire IL1_D3_LR1_D3_read_en;
wire [35:0] IL1_D3_LR1_D3;
//wire IL1_D3_LR1_D3_empty;
InputLink  IL1_D3(
.data_in1(input_link1_reg1),
.data_in2(input_link1_reg2),
.read_en(IL1_D3_LR1_D3_read_en),
.data_out(IL1_D3_LR1_D3),
.empty(IL1_D3_LR1_D3_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire IL2_D3_LR2_D3_read_en;
wire [35:0] IL2_D3_LR2_D3;
//wire IL2_D3_LR2_D3_empty;
InputLink  IL2_D3(
.data_in1(input_link2_reg1),
.data_in2(input_link2_reg2),
.read_en(IL2_D3_LR2_D3_read_en),
.data_out(IL2_D3_LR2_D3),
.empty(IL2_D3_LR2_D3_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire IL3_D3_LR3_D3_read_en;
wire [35:0] IL3_D3_LR3_D3;
//wire IL3_D3_LR3_D3_empty;
InputLink  IL3_D3(
.data_in1(input_link3_reg1),
.data_in2(input_link3_reg2),
.read_en(IL3_D3_LR3_D3_read_en),
.data_out(IL3_D3_LR3_D3),
.empty(IL3_D3_LR3_D3_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire IL1_D4_LR1_D4_read_en;
wire [35:0] IL1_D4_LR1_D4;
//wire IL1_D4_LR1_D4_empty;
InputLink  IL1_D4(
.data_in1(input_link4_reg1),
.data_in2(input_link4_reg2),
.read_en(IL1_D4_LR1_D4_read_en),
.data_out(IL1_D4_LR1_D4),
.empty(IL1_D4_LR1_D4_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire IL2_D4_LR2_D4_read_en;
wire [35:0] IL2_D4_LR2_D4;
//wire IL2_D4_LR2_D4_empty;
InputLink  IL2_D4(
.data_in1(input_link5_reg1),
.data_in2(input_link5_reg2),
.read_en(IL2_D4_LR2_D4_read_en),
.data_out(IL2_D4_LR2_D4),
.empty(IL2_D4_LR2_D4_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire IL3_D4_LR3_D4_read_en;
wire [35:0] IL3_D4_LR3_D4;
//wire IL3_D4_LR3_D4_empty;
InputLink  IL3_D4(
.data_in1(input_link6_reg1),
.data_in2(input_link6_reg2),
.read_en(IL3_D4_LR3_D4_read_en),
.data_out(IL3_D4_LR3_D4),
.empty(IL3_D4_LR3_D4_empty),
.start(),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D3_SL1_L1D3;
wire LR1_D3_SL1_L1D3_wr_en;
wire [5:0] SL1_L1D3_VMR_L1D3_number;
wire [8:0] SL1_L1D3_VMR_L1D3_read_add;
wire [35:0] SL1_L1D3_VMR_L1D3;
StubsByLayer  SL1_L1D3(
.data_in(LR1_D3_SL1_L1D3),
.enable(LR1_D3_SL1_L1D3_wr_en),
.number_out(SL1_L1D3_VMR_L1D3_number),
.read_add(SL1_L1D3_VMR_L1D3_read_add),
.data_out(SL1_L1D3_VMR_L1D3),
.start(LR1_D3_start),
.done(SL1_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D3_SL2_L1D3;
wire LR2_D3_SL2_L1D3_wr_en;
wire [5:0] SL2_L1D3_VMR_L1D3_number;
wire [8:0] SL2_L1D3_VMR_L1D3_read_add;
wire [35:0] SL2_L1D3_VMR_L1D3;
StubsByLayer  SL2_L1D3(
.data_in(LR2_D3_SL2_L1D3),
.enable(LR2_D3_SL2_L1D3_wr_en),
.number_out(SL2_L1D3_VMR_L1D3_number),
.read_add(SL2_L1D3_VMR_L1D3_read_add),
.data_out(SL2_L1D3_VMR_L1D3),
.start(LR2_D3_start),
.done(SL2_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D3_SL3_L1D3;
wire LR3_D3_SL3_L1D3_wr_en;
wire [5:0] SL3_L1D3_VMR_L1D3_number;
wire [8:0] SL3_L1D3_VMR_L1D3_read_add;
wire [35:0] SL3_L1D3_VMR_L1D3;
StubsByLayer  SL3_L1D3(
.data_in(LR3_D3_SL3_L1D3),
.enable(LR3_D3_SL3_L1D3_wr_en),
.number_out(SL3_L1D3_VMR_L1D3_number),
.read_add(SL3_L1D3_VMR_L1D3_read_add),
.data_out(SL3_L1D3_VMR_L1D3),
.start(LR3_D3_start),
.done(SL3_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D4_SL1_L1D4;
wire LR1_D4_SL1_L1D4_wr_en;
wire [5:0] SL1_L1D4_VMR_L1D4_number;
wire [8:0] SL1_L1D4_VMR_L1D4_read_add;
wire [35:0] SL1_L1D4_VMR_L1D4;
StubsByLayer  SL1_L1D4(
.data_in(LR1_D4_SL1_L1D4),
.enable(LR1_D4_SL1_L1D4_wr_en),
.number_out(SL1_L1D4_VMR_L1D4_number),
.read_add(SL1_L1D4_VMR_L1D4_read_add),
.data_out(SL1_L1D4_VMR_L1D4),
.start(LR1_D4_start),
.done(SL1_L1D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D4_SL2_L1D4;
wire LR2_D4_SL2_L1D4_wr_en;
wire [5:0] SL2_L1D4_VMR_L1D4_number;
wire [8:0] SL2_L1D4_VMR_L1D4_read_add;
wire [35:0] SL2_L1D4_VMR_L1D4;
StubsByLayer  SL2_L1D4(
.data_in(LR2_D4_SL2_L1D4),
.enable(LR2_D4_SL2_L1D4_wr_en),
.number_out(SL2_L1D4_VMR_L1D4_number),
.read_add(SL2_L1D4_VMR_L1D4_read_add),
.data_out(SL2_L1D4_VMR_L1D4),
.start(LR2_D4_start),
.done(SL2_L1D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D4_SL3_L1D4;
wire LR3_D4_SL3_L1D4_wr_en;
wire [5:0] SL3_L1D4_VMR_L1D4_number;
wire [8:0] SL3_L1D4_VMR_L1D4_read_add;
wire [35:0] SL3_L1D4_VMR_L1D4;
StubsByLayer  SL3_L1D4(
.data_in(LR3_D4_SL3_L1D4),
.enable(LR3_D4_SL3_L1D4_wr_en),
.number_out(SL3_L1D4_VMR_L1D4_number),
.read_add(SL3_L1D4_VMR_L1D4_read_add),
.data_out(SL3_L1D4_VMR_L1D4),
.start(LR3_D4_start),
.done(SL3_L1D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D3_SL1_L2D3;
wire LR1_D3_SL1_L2D3_wr_en;
wire [5:0] SL1_L2D3_VMR_L2D3_number;
wire [8:0] SL1_L2D3_VMR_L2D3_read_add;
wire [35:0] SL1_L2D3_VMR_L2D3;
StubsByLayer  SL1_L2D3(
.data_in(LR1_D3_SL1_L2D3),
.enable(LR1_D3_SL1_L2D3_wr_en),
.number_out(SL1_L2D3_VMR_L2D3_number),
.read_add(SL1_L2D3_VMR_L2D3_read_add),
.data_out(SL1_L2D3_VMR_L2D3),
.start(LR1_D3_start),
.done(SL1_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D3_SL2_L2D3;
wire LR2_D3_SL2_L2D3_wr_en;
wire [5:0] SL2_L2D3_VMR_L2D3_number;
wire [8:0] SL2_L2D3_VMR_L2D3_read_add;
wire [35:0] SL2_L2D3_VMR_L2D3;
StubsByLayer  SL2_L2D3(
.data_in(LR2_D3_SL2_L2D3),
.enable(LR2_D3_SL2_L2D3_wr_en),
.number_out(SL2_L2D3_VMR_L2D3_number),
.read_add(SL2_L2D3_VMR_L2D3_read_add),
.data_out(SL2_L2D3_VMR_L2D3),
.start(LR2_D3_start),
.done(SL2_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D3_SL3_L2D3;
wire LR3_D3_SL3_L2D3_wr_en;
wire [5:0] SL3_L2D3_VMR_L2D3_number;
wire [8:0] SL3_L2D3_VMR_L2D3_read_add;
wire [35:0] SL3_L2D3_VMR_L2D3;
StubsByLayer  SL3_L2D3(
.data_in(LR3_D3_SL3_L2D3),
.enable(LR3_D3_SL3_L2D3_wr_en),
.number_out(SL3_L2D3_VMR_L2D3_number),
.read_add(SL3_L2D3_VMR_L2D3_read_add),
.data_out(SL3_L2D3_VMR_L2D3),
.start(LR3_D3_start),
.done(SL3_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D4_SL1_L2D4;
wire LR1_D4_SL1_L2D4_wr_en;
wire [5:0] SL1_L2D4_VMR_L2D4_number;
wire [8:0] SL1_L2D4_VMR_L2D4_read_add;
wire [35:0] SL1_L2D4_VMR_L2D4;
StubsByLayer  SL1_L2D4(
.data_in(LR1_D4_SL1_L2D4),
.enable(LR1_D4_SL1_L2D4_wr_en),
.number_out(SL1_L2D4_VMR_L2D4_number),
.read_add(SL1_L2D4_VMR_L2D4_read_add),
.data_out(SL1_L2D4_VMR_L2D4),
.start(LR1_D4_start),
.done(SL1_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D4_SL2_L2D4;
wire LR2_D4_SL2_L2D4_wr_en;
wire [5:0] SL2_L2D4_VMR_L2D4_number;
wire [8:0] SL2_L2D4_VMR_L2D4_read_add;
wire [35:0] SL2_L2D4_VMR_L2D4;
StubsByLayer  SL2_L2D4(
.data_in(LR2_D4_SL2_L2D4),
.enable(LR2_D4_SL2_L2D4_wr_en),
.number_out(SL2_L2D4_VMR_L2D4_number),
.read_add(SL2_L2D4_VMR_L2D4_read_add),
.data_out(SL2_L2D4_VMR_L2D4),
.start(LR2_D4_start),
.done(SL2_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D4_SL3_L2D4;
wire LR3_D4_SL3_L2D4_wr_en;
wire [5:0] SL3_L2D4_VMR_L2D4_number;
wire [8:0] SL3_L2D4_VMR_L2D4_read_add;
wire [35:0] SL3_L2D4_VMR_L2D4;
StubsByLayer  SL3_L2D4(
.data_in(LR3_D4_SL3_L2D4),
.enable(LR3_D4_SL3_L2D4_wr_en),
.number_out(SL3_L2D4_VMR_L2D4_number),
.read_add(SL3_L2D4_VMR_L2D4_read_add),
.data_out(SL3_L2D4_VMR_L2D4),
.start(LR3_D4_start),
.done(SL3_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D3_SL1_L3D3;
wire LR1_D3_SL1_L3D3_wr_en;
wire [5:0] SL1_L3D3_VMR_L3D3_number;
wire [8:0] SL1_L3D3_VMR_L3D3_read_add;
wire [35:0] SL1_L3D3_VMR_L3D3;
StubsByLayer  SL1_L3D3(
.data_in(LR1_D3_SL1_L3D3),
.enable(LR1_D3_SL1_L3D3_wr_en),
.number_out(SL1_L3D3_VMR_L3D3_number),
.read_add(SL1_L3D3_VMR_L3D3_read_add),
.data_out(SL1_L3D3_VMR_L3D3),
.start(LR1_D3_start),
.done(SL1_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D3_SL2_L3D3;
wire LR2_D3_SL2_L3D3_wr_en;
wire [5:0] SL2_L3D3_VMR_L3D3_number;
wire [8:0] SL2_L3D3_VMR_L3D3_read_add;
wire [35:0] SL2_L3D3_VMR_L3D3;
StubsByLayer  SL2_L3D3(
.data_in(LR2_D3_SL2_L3D3),
.enable(LR2_D3_SL2_L3D3_wr_en),
.number_out(SL2_L3D3_VMR_L3D3_number),
.read_add(SL2_L3D3_VMR_L3D3_read_add),
.data_out(SL2_L3D3_VMR_L3D3),
.start(LR2_D3_start),
.done(SL2_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D3_SL3_L3D3;
wire LR3_D3_SL3_L3D3_wr_en;
wire [5:0] SL3_L3D3_VMR_L3D3_number;
wire [8:0] SL3_L3D3_VMR_L3D3_read_add;
wire [35:0] SL3_L3D3_VMR_L3D3;
StubsByLayer  SL3_L3D3(
.data_in(LR3_D3_SL3_L3D3),
.enable(LR3_D3_SL3_L3D3_wr_en),
.number_out(SL3_L3D3_VMR_L3D3_number),
.read_add(SL3_L3D3_VMR_L3D3_read_add),
.data_out(SL3_L3D3_VMR_L3D3),
.start(LR3_D3_start),
.done(SL3_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D4_SL1_L3D4;
wire LR1_D4_SL1_L3D4_wr_en;
wire [5:0] SL1_L3D4_VMR_L3D4_number;
wire [8:0] SL1_L3D4_VMR_L3D4_read_add;
wire [35:0] SL1_L3D4_VMR_L3D4;
StubsByLayer  SL1_L3D4(
.data_in(LR1_D4_SL1_L3D4),
.enable(LR1_D4_SL1_L3D4_wr_en),
.number_out(SL1_L3D4_VMR_L3D4_number),
.read_add(SL1_L3D4_VMR_L3D4_read_add),
.data_out(SL1_L3D4_VMR_L3D4),
.start(LR1_D4_start),
.done(SL1_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D4_SL2_L3D4;
wire LR2_D4_SL2_L3D4_wr_en;
wire [5:0] SL2_L3D4_VMR_L3D4_number;
wire [8:0] SL2_L3D4_VMR_L3D4_read_add;
wire [35:0] SL2_L3D4_VMR_L3D4;
StubsByLayer  SL2_L3D4(
.data_in(LR2_D4_SL2_L3D4),
.enable(LR2_D4_SL2_L3D4_wr_en),
.number_out(SL2_L3D4_VMR_L3D4_number),
.read_add(SL2_L3D4_VMR_L3D4_read_add),
.data_out(SL2_L3D4_VMR_L3D4),
.start(LR2_D4_start),
.done(SL2_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D4_SL3_L3D4;
wire LR3_D4_SL3_L3D4_wr_en;
wire [5:0] SL3_L3D4_VMR_L3D4_number;
wire [8:0] SL3_L3D4_VMR_L3D4_read_add;
wire [35:0] SL3_L3D4_VMR_L3D4;
StubsByLayer  SL3_L3D4(
.data_in(LR3_D4_SL3_L3D4),
.enable(LR3_D4_SL3_L3D4_wr_en),
.number_out(SL3_L3D4_VMR_L3D4_number),
.read_add(SL3_L3D4_VMR_L3D4_read_add),
.data_out(SL3_L3D4_VMR_L3D4),
.start(LR3_D4_start),
.done(SL3_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D3_SL1_L4D3;
wire LR1_D3_SL1_L4D3_wr_en;
wire [5:0] SL1_L4D3_VMR_L4D3_number;
wire [8:0] SL1_L4D3_VMR_L4D3_read_add;
wire [35:0] SL1_L4D3_VMR_L4D3;
StubsByLayer  SL1_L4D3(
.data_in(LR1_D3_SL1_L4D3),
.enable(LR1_D3_SL1_L4D3_wr_en),
.number_out(SL1_L4D3_VMR_L4D3_number),
.read_add(SL1_L4D3_VMR_L4D3_read_add),
.data_out(SL1_L4D3_VMR_L4D3),
.start(LR1_D3_start),
.done(SL1_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D3_SL2_L4D3;
wire LR2_D3_SL2_L4D3_wr_en;
wire [5:0] SL2_L4D3_VMR_L4D3_number;
wire [8:0] SL2_L4D3_VMR_L4D3_read_add;
wire [35:0] SL2_L4D3_VMR_L4D3;
StubsByLayer  SL2_L4D3(
.data_in(LR2_D3_SL2_L4D3),
.enable(LR2_D3_SL2_L4D3_wr_en),
.number_out(SL2_L4D3_VMR_L4D3_number),
.read_add(SL2_L4D3_VMR_L4D3_read_add),
.data_out(SL2_L4D3_VMR_L4D3),
.start(LR2_D3_start),
.done(SL2_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D3_SL3_L4D3;
wire LR3_D3_SL3_L4D3_wr_en;
wire [5:0] SL3_L4D3_VMR_L4D3_number;
wire [8:0] SL3_L4D3_VMR_L4D3_read_add;
wire [35:0] SL3_L4D3_VMR_L4D3;
StubsByLayer  SL3_L4D3(
.data_in(LR3_D3_SL3_L4D3),
.enable(LR3_D3_SL3_L4D3_wr_en),
.number_out(SL3_L4D3_VMR_L4D3_number),
.read_add(SL3_L4D3_VMR_L4D3_read_add),
.data_out(SL3_L4D3_VMR_L4D3),
.start(LR3_D3_start),
.done(SL3_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D4_SL1_L4D4;
wire LR1_D4_SL1_L4D4_wr_en;
wire [5:0] SL1_L4D4_VMR_L4D4_number;
wire [8:0] SL1_L4D4_VMR_L4D4_read_add;
wire [35:0] SL1_L4D4_VMR_L4D4;
StubsByLayer  SL1_L4D4(
.data_in(LR1_D4_SL1_L4D4),
.enable(LR1_D4_SL1_L4D4_wr_en),
.number_out(SL1_L4D4_VMR_L4D4_number),
.read_add(SL1_L4D4_VMR_L4D4_read_add),
.data_out(SL1_L4D4_VMR_L4D4),
.start(LR1_D4_start),
.done(SL1_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D4_SL2_L4D4;
wire LR2_D4_SL2_L4D4_wr_en;
wire [5:0] SL2_L4D4_VMR_L4D4_number;
wire [8:0] SL2_L4D4_VMR_L4D4_read_add;
wire [35:0] SL2_L4D4_VMR_L4D4;
StubsByLayer  SL2_L4D4(
.data_in(LR2_D4_SL2_L4D4),
.enable(LR2_D4_SL2_L4D4_wr_en),
.number_out(SL2_L4D4_VMR_L4D4_number),
.read_add(SL2_L4D4_VMR_L4D4_read_add),
.data_out(SL2_L4D4_VMR_L4D4),
.start(LR2_D4_start),
.done(SL2_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D4_SL3_L4D4;
wire LR3_D4_SL3_L4D4_wr_en;
wire [5:0] SL3_L4D4_VMR_L4D4_number;
wire [8:0] SL3_L4D4_VMR_L4D4_read_add;
wire [35:0] SL3_L4D4_VMR_L4D4;
StubsByLayer  SL3_L4D4(
.data_in(LR3_D4_SL3_L4D4),
.enable(LR3_D4_SL3_L4D4_wr_en),
.number_out(SL3_L4D4_VMR_L4D4_number),
.read_add(SL3_L4D4_VMR_L4D4_read_add),
.data_out(SL3_L4D4_VMR_L4D4),
.start(LR3_D4_start),
.done(SL3_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D3_SL1_L5D3;
wire LR1_D3_SL1_L5D3_wr_en;
wire [5:0] SL1_L5D3_VMR_L5D3_number;
wire [8:0] SL1_L5D3_VMR_L5D3_read_add;
wire [35:0] SL1_L5D3_VMR_L5D3;
StubsByLayer  SL1_L5D3(
.data_in(LR1_D3_SL1_L5D3),
.enable(LR1_D3_SL1_L5D3_wr_en),
.number_out(SL1_L5D3_VMR_L5D3_number),
.read_add(SL1_L5D3_VMR_L5D3_read_add),
.data_out(SL1_L5D3_VMR_L5D3),
.start(LR1_D3_start),
.done(SL1_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D3_SL2_L5D3;
wire LR2_D3_SL2_L5D3_wr_en;
wire [5:0] SL2_L5D3_VMR_L5D3_number;
wire [8:0] SL2_L5D3_VMR_L5D3_read_add;
wire [35:0] SL2_L5D3_VMR_L5D3;
StubsByLayer  SL2_L5D3(
.data_in(LR2_D3_SL2_L5D3),
.enable(LR2_D3_SL2_L5D3_wr_en),
.number_out(SL2_L5D3_VMR_L5D3_number),
.read_add(SL2_L5D3_VMR_L5D3_read_add),
.data_out(SL2_L5D3_VMR_L5D3),
.start(LR2_D3_start),
.done(SL2_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D3_SL3_L5D3;
wire LR3_D3_SL3_L5D3_wr_en;
wire [5:0] SL3_L5D3_VMR_L5D3_number;
wire [8:0] SL3_L5D3_VMR_L5D3_read_add;
wire [35:0] SL3_L5D3_VMR_L5D3;
StubsByLayer  SL3_L5D3(
.data_in(LR3_D3_SL3_L5D3),
.enable(LR3_D3_SL3_L5D3_wr_en),
.number_out(SL3_L5D3_VMR_L5D3_number),
.read_add(SL3_L5D3_VMR_L5D3_read_add),
.data_out(SL3_L5D3_VMR_L5D3),
.start(LR3_D3_start),
.done(SL3_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D4_SL1_L5D4;
wire LR1_D4_SL1_L5D4_wr_en;
wire [5:0] SL1_L5D4_VMR_L5D4_number;
wire [8:0] SL1_L5D4_VMR_L5D4_read_add;
wire [35:0] SL1_L5D4_VMR_L5D4;
StubsByLayer  SL1_L5D4(
.data_in(LR1_D4_SL1_L5D4),
.enable(LR1_D4_SL1_L5D4_wr_en),
.number_out(SL1_L5D4_VMR_L5D4_number),
.read_add(SL1_L5D4_VMR_L5D4_read_add),
.data_out(SL1_L5D4_VMR_L5D4),
.start(LR1_D4_start),
.done(SL1_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D4_SL2_L5D4;
wire LR2_D4_SL2_L5D4_wr_en;
wire [5:0] SL2_L5D4_VMR_L5D4_number;
wire [8:0] SL2_L5D4_VMR_L5D4_read_add;
wire [35:0] SL2_L5D4_VMR_L5D4;
StubsByLayer  SL2_L5D4(
.data_in(LR2_D4_SL2_L5D4),
.enable(LR2_D4_SL2_L5D4_wr_en),
.number_out(SL2_L5D4_VMR_L5D4_number),
.read_add(SL2_L5D4_VMR_L5D4_read_add),
.data_out(SL2_L5D4_VMR_L5D4),
.start(LR2_D4_start),
.done(SL2_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D4_SL3_L5D4;
wire LR3_D4_SL3_L5D4_wr_en;
wire [5:0] SL3_L5D4_VMR_L5D4_number;
wire [8:0] SL3_L5D4_VMR_L5D4_read_add;
wire [35:0] SL3_L5D4_VMR_L5D4;
StubsByLayer  SL3_L5D4(
.data_in(LR3_D4_SL3_L5D4),
.enable(LR3_D4_SL3_L5D4_wr_en),
.number_out(SL3_L5D4_VMR_L5D4_number),
.read_add(SL3_L5D4_VMR_L5D4_read_add),
.data_out(SL3_L5D4_VMR_L5D4),
.start(LR3_D4_start),
.done(SL3_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D3_SL1_L6D3;
wire LR1_D3_SL1_L6D3_wr_en;
wire [5:0] SL1_L6D3_VMR_L6D3_number;
wire [8:0] SL1_L6D3_VMR_L6D3_read_add;
wire [35:0] SL1_L6D3_VMR_L6D3;
StubsByLayer  SL1_L6D3(
.data_in(LR1_D3_SL1_L6D3),
.enable(LR1_D3_SL1_L6D3_wr_en),
.number_out(SL1_L6D3_VMR_L6D3_number),
.read_add(SL1_L6D3_VMR_L6D3_read_add),
.data_out(SL1_L6D3_VMR_L6D3),
.start(LR1_D3_start),
.done(SL1_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D3_SL2_L6D3;
wire LR2_D3_SL2_L6D3_wr_en;
wire [5:0] SL2_L6D3_VMR_L6D3_number;
wire [8:0] SL2_L6D3_VMR_L6D3_read_add;
wire [35:0] SL2_L6D3_VMR_L6D3;
StubsByLayer  SL2_L6D3(
.data_in(LR2_D3_SL2_L6D3),
.enable(LR2_D3_SL2_L6D3_wr_en),
.number_out(SL2_L6D3_VMR_L6D3_number),
.read_add(SL2_L6D3_VMR_L6D3_read_add),
.data_out(SL2_L6D3_VMR_L6D3),
.start(LR2_D3_start),
.done(SL2_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D3_SL3_L6D3;
wire LR3_D3_SL3_L6D3_wr_en;
wire [5:0] SL3_L6D3_VMR_L6D3_number;
wire [8:0] SL3_L6D3_VMR_L6D3_read_add;
wire [35:0] SL3_L6D3_VMR_L6D3;
StubsByLayer  SL3_L6D3(
.data_in(LR3_D3_SL3_L6D3),
.enable(LR3_D3_SL3_L6D3_wr_en),
.number_out(SL3_L6D3_VMR_L6D3_number),
.read_add(SL3_L6D3_VMR_L6D3_read_add),
.data_out(SL3_L6D3_VMR_L6D3),
.start(LR3_D3_start),
.done(SL3_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR1_D4_SL1_L6D4;
wire LR1_D4_SL1_L6D4_wr_en;
wire [5:0] SL1_L6D4_VMR_L6D4_number;
wire [8:0] SL1_L6D4_VMR_L6D4_read_add;
wire [35:0] SL1_L6D4_VMR_L6D4;
StubsByLayer  SL1_L6D4(
.data_in(LR1_D4_SL1_L6D4),
.enable(LR1_D4_SL1_L6D4_wr_en),
.number_out(SL1_L6D4_VMR_L6D4_number),
.read_add(SL1_L6D4_VMR_L6D4_read_add),
.data_out(SL1_L6D4_VMR_L6D4),
.start(LR1_D4_start),
.done(SL1_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR2_D4_SL2_L6D4;
wire LR2_D4_SL2_L6D4_wr_en;
wire [5:0] SL2_L6D4_VMR_L6D4_number;
wire [8:0] SL2_L6D4_VMR_L6D4_read_add;
wire [35:0] SL2_L6D4_VMR_L6D4;
StubsByLayer  SL2_L6D4(
.data_in(LR2_D4_SL2_L6D4),
.enable(LR2_D4_SL2_L6D4_wr_en),
.number_out(SL2_L6D4_VMR_L6D4_number),
.read_add(SL2_L6D4_VMR_L6D4_read_add),
.data_out(SL2_L6D4_VMR_L6D4),
.start(LR2_D4_start),
.done(SL2_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] LR3_D4_SL3_L6D4;
wire LR3_D4_SL3_L6D4_wr_en;
wire [5:0] SL3_L6D4_VMR_L6D4_number;
wire [8:0] SL3_L6D4_VMR_L6D4_read_add;
wire [35:0] SL3_L6D4_VMR_L6D4;
StubsByLayer  SL3_L6D4(
.data_in(LR3_D4_SL3_L6D4),
.enable(LR3_D4_SL3_L6D4_wr_en),
.number_out(SL3_L6D4_VMR_L6D4_number),
.read_add(SL3_L6D4_VMR_L6D4_read_add),
.data_out(SL3_L6D4_VMR_L6D4),
.start(LR3_D4_start),
.done(SL3_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X1n1;
wire VMR_L1D3_VMS_L1D3PHI1X1n1_wr_en;
wire [5:0] VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_number;
wire [10:0] VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_read_add;
wire [18:0] VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1;
VMStubs #("Tracklet") VMS_L1D3PHI1X1n1(
.data_in(VMR_L1D3_VMS_L1D3PHI1X1n1),
.enable(VMR_L1D3_VMS_L1D3PHI1X1n1_wr_en),
.number_out(VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_number),
.read_add(VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_read_add),
.data_out(VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI1X1n1;
wire VMR_L2D3_VMS_L2D3PHI1X1n1_wr_en;
wire [5:0] VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_number;
wire [10:0] VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_read_add;
wire [18:0] VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1;
VMStubs #("Tracklet") VMS_L2D3PHI1X1n1(
.data_in(VMR_L2D3_VMS_L2D3PHI1X1n1),
.enable(VMR_L2D3_VMS_L2D3PHI1X1n1_wr_en),
.number_out(VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_number),
.read_add(VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_read_add),
.data_out(VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X1n2;
wire VMR_L1D3_VMS_L1D3PHI1X1n2_wr_en;
wire [5:0] VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1_number;
wire [10:0] VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1_read_add;
wire [18:0] VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1;
VMStubs #("Tracklet") VMS_L1D3PHI1X1n2(
.data_in(VMR_L1D3_VMS_L1D3PHI1X1n2),
.enable(VMR_L1D3_VMS_L1D3PHI1X1n2_wr_en),
.number_out(VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1_number),
.read_add(VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1_read_add),
.data_out(VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X1n1;
wire VMR_L2D3_VMS_L2D3PHI2X1n1_wr_en;
wire [5:0] VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1_number;
wire [10:0] VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1_read_add;
wire [18:0] VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1;
VMStubs #("Tracklet") VMS_L2D3PHI2X1n1(
.data_in(VMR_L2D3_VMS_L2D3PHI2X1n1),
.enable(VMR_L2D3_VMS_L2D3PHI2X1n1_wr_en),
.number_out(VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1_number),
.read_add(VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1_read_add),
.data_out(VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X1n1;
wire VMR_L1D3_VMS_L1D3PHI2X1n1_wr_en;
wire [5:0] VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1_number;
wire [10:0] VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1_read_add;
wire [18:0] VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1;
VMStubs #("Tracklet") VMS_L1D3PHI2X1n1(
.data_in(VMR_L1D3_VMS_L1D3PHI2X1n1),
.enable(VMR_L1D3_VMS_L1D3PHI2X1n1_wr_en),
.number_out(VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1_number),
.read_add(VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1_read_add),
.data_out(VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X1n2;
wire VMR_L2D3_VMS_L2D3PHI2X1n2_wr_en;
wire [5:0] VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1_number;
wire [10:0] VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1_read_add;
wire [18:0] VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1;
VMStubs #("Tracklet") VMS_L2D3PHI2X1n2(
.data_in(VMR_L2D3_VMS_L2D3PHI2X1n2),
.enable(VMR_L2D3_VMS_L2D3PHI2X1n2_wr_en),
.number_out(VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1_number),
.read_add(VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1_read_add),
.data_out(VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X1n2;
wire VMR_L1D3_VMS_L1D3PHI2X1n2_wr_en;
wire [5:0] VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1_number;
wire [10:0] VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1_read_add;
wire [18:0] VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1;
VMStubs #("Tracklet") VMS_L1D3PHI2X1n2(
.data_in(VMR_L1D3_VMS_L1D3PHI2X1n2),
.enable(VMR_L1D3_VMS_L1D3PHI2X1n2_wr_en),
.number_out(VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1_number),
.read_add(VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1_read_add),
.data_out(VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X1n1;
wire VMR_L2D3_VMS_L2D3PHI3X1n1_wr_en;
wire [5:0] VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1_number;
wire [10:0] VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1_read_add;
wire [18:0] VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1;
VMStubs #("Tracklet") VMS_L2D3PHI3X1n1(
.data_in(VMR_L2D3_VMS_L2D3PHI3X1n1),
.enable(VMR_L2D3_VMS_L2D3PHI3X1n1_wr_en),
.number_out(VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1_number),
.read_add(VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1_read_add),
.data_out(VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X1n1;
wire VMR_L1D3_VMS_L1D3PHI3X1n1_wr_en;
wire [5:0] VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1_number;
wire [10:0] VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1_read_add;
wire [18:0] VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1;
VMStubs #("Tracklet") VMS_L1D3PHI3X1n1(
.data_in(VMR_L1D3_VMS_L1D3PHI3X1n1),
.enable(VMR_L1D3_VMS_L1D3PHI3X1n1_wr_en),
.number_out(VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1_number),
.read_add(VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1_read_add),
.data_out(VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X1n2;
wire VMR_L2D3_VMS_L2D3PHI3X1n2_wr_en;
wire [5:0] VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1_number;
wire [10:0] VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1_read_add;
wire [18:0] VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1;
VMStubs #("Tracklet") VMS_L2D3PHI3X1n2(
.data_in(VMR_L2D3_VMS_L2D3PHI3X1n2),
.enable(VMR_L2D3_VMS_L2D3PHI3X1n2_wr_en),
.number_out(VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1_number),
.read_add(VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1_read_add),
.data_out(VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X1n2;
wire VMR_L1D3_VMS_L1D3PHI3X1n2_wr_en;
wire [5:0] VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1_number;
wire [10:0] VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1_read_add;
wire [18:0] VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1;
VMStubs #("Tracklet") VMS_L1D3PHI3X1n2(
.data_in(VMR_L1D3_VMS_L1D3PHI3X1n2),
.enable(VMR_L1D3_VMS_L1D3PHI3X1n2_wr_en),
.number_out(VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1_number),
.read_add(VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1_read_add),
.data_out(VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI4X1n1;
wire VMR_L2D3_VMS_L2D3PHI4X1n1_wr_en;
wire [5:0] VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1_number;
wire [10:0] VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1_read_add;
wire [18:0] VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1;
VMStubs #("Tracklet") VMS_L2D3PHI4X1n1(
.data_in(VMR_L2D3_VMS_L2D3PHI4X1n1),
.enable(VMR_L2D3_VMS_L2D3PHI4X1n1_wr_en),
.number_out(VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1_number),
.read_add(VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1_read_add),
.data_out(VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X1n3;
wire VMR_L1D3_VMS_L1D3PHI1X1n3_wr_en;
wire [5:0] VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2_number;
wire [10:0] VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2_read_add;
wire [18:0] VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2;
VMStubs #("Tracklet") VMS_L1D3PHI1X1n3(
.data_in(VMR_L1D3_VMS_L1D3PHI1X1n3),
.enable(VMR_L1D3_VMS_L1D3PHI1X1n3_wr_en),
.number_out(VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2_number),
.read_add(VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2_read_add),
.data_out(VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI1X2n1;
wire VMR_L2D3_VMS_L2D3PHI1X2n1_wr_en;
wire [5:0] VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2_number;
wire [10:0] VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2_read_add;
wire [18:0] VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2;
VMStubs #("Tracklet") VMS_L2D3PHI1X2n1(
.data_in(VMR_L2D3_VMS_L2D3PHI1X2n1),
.enable(VMR_L2D3_VMS_L2D3PHI1X2n1_wr_en),
.number_out(VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2_number),
.read_add(VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2_read_add),
.data_out(VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X1n4;
wire VMR_L1D3_VMS_L1D3PHI1X1n4_wr_en;
wire [5:0] VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2_number;
wire [10:0] VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2_read_add;
wire [18:0] VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2;
VMStubs #("Tracklet") VMS_L1D3PHI1X1n4(
.data_in(VMR_L1D3_VMS_L1D3PHI1X1n4),
.enable(VMR_L1D3_VMS_L1D3PHI1X1n4_wr_en),
.number_out(VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2_number),
.read_add(VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2_read_add),
.data_out(VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X2n1;
wire VMR_L2D3_VMS_L2D3PHI2X2n1_wr_en;
wire [5:0] VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2_number;
wire [10:0] VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2_read_add;
wire [18:0] VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2;
VMStubs #("Tracklet") VMS_L2D3PHI2X2n1(
.data_in(VMR_L2D3_VMS_L2D3PHI2X2n1),
.enable(VMR_L2D3_VMS_L2D3PHI2X2n1_wr_en),
.number_out(VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2_number),
.read_add(VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2_read_add),
.data_out(VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X1n3;
wire VMR_L1D3_VMS_L1D3PHI2X1n3_wr_en;
wire [5:0] VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2_number;
wire [10:0] VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2_read_add;
wire [18:0] VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2;
VMStubs #("Tracklet") VMS_L1D3PHI2X1n3(
.data_in(VMR_L1D3_VMS_L1D3PHI2X1n3),
.enable(VMR_L1D3_VMS_L1D3PHI2X1n3_wr_en),
.number_out(VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2_number),
.read_add(VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2_read_add),
.data_out(VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X2n2;
wire VMR_L2D3_VMS_L2D3PHI2X2n2_wr_en;
wire [5:0] VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2_number;
wire [10:0] VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2_read_add;
wire [18:0] VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2;
VMStubs #("Tracklet") VMS_L2D3PHI2X2n2(
.data_in(VMR_L2D3_VMS_L2D3PHI2X2n2),
.enable(VMR_L2D3_VMS_L2D3PHI2X2n2_wr_en),
.number_out(VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2_number),
.read_add(VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2_read_add),
.data_out(VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X1n4;
wire VMR_L1D3_VMS_L1D3PHI2X1n4_wr_en;
wire [5:0] VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2_number;
wire [10:0] VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2_read_add;
wire [18:0] VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2;
VMStubs #("Tracklet") VMS_L1D3PHI2X1n4(
.data_in(VMR_L1D3_VMS_L1D3PHI2X1n4),
.enable(VMR_L1D3_VMS_L1D3PHI2X1n4_wr_en),
.number_out(VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2_number),
.read_add(VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2_read_add),
.data_out(VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X2n1;
wire VMR_L2D3_VMS_L2D3PHI3X2n1_wr_en;
wire [5:0] VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2_number;
wire [10:0] VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2_read_add;
wire [18:0] VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2;
VMStubs #("Tracklet") VMS_L2D3PHI3X2n1(
.data_in(VMR_L2D3_VMS_L2D3PHI3X2n1),
.enable(VMR_L2D3_VMS_L2D3PHI3X2n1_wr_en),
.number_out(VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2_number),
.read_add(VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2_read_add),
.data_out(VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X1n3;
wire VMR_L1D3_VMS_L1D3PHI3X1n3_wr_en;
wire [5:0] VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2_number;
wire [10:0] VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2_read_add;
wire [18:0] VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2;
VMStubs #("Tracklet") VMS_L1D3PHI3X1n3(
.data_in(VMR_L1D3_VMS_L1D3PHI3X1n3),
.enable(VMR_L1D3_VMS_L1D3PHI3X1n3_wr_en),
.number_out(VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2_number),
.read_add(VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2_read_add),
.data_out(VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X2n2;
wire VMR_L2D3_VMS_L2D3PHI3X2n2_wr_en;
wire [5:0] VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2_number;
wire [10:0] VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2_read_add;
wire [18:0] VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2;
VMStubs #("Tracklet") VMS_L2D3PHI3X2n2(
.data_in(VMR_L2D3_VMS_L2D3PHI3X2n2),
.enable(VMR_L2D3_VMS_L2D3PHI3X2n2_wr_en),
.number_out(VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2_number),
.read_add(VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2_read_add),
.data_out(VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X1n4;
wire VMR_L1D3_VMS_L1D3PHI3X1n4_wr_en;
wire [5:0] VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2_number;
wire [10:0] VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2_read_add;
wire [18:0] VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2;
VMStubs #("Tracklet") VMS_L1D3PHI3X1n4(
.data_in(VMR_L1D3_VMS_L1D3PHI3X1n4),
.enable(VMR_L1D3_VMS_L1D3PHI3X1n4_wr_en),
.number_out(VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2_number),
.read_add(VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2_read_add),
.data_out(VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI4X2n1;
wire VMR_L2D3_VMS_L2D3PHI4X2n1_wr_en;
wire [5:0] VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2_number;
wire [10:0] VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2_read_add;
wire [18:0] VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2;
VMStubs #("Tracklet") VMS_L2D3PHI4X2n1(
.data_in(VMR_L2D3_VMS_L2D3PHI4X2n1),
.enable(VMR_L2D3_VMS_L2D3PHI4X2n1_wr_en),
.number_out(VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2_number),
.read_add(VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2_read_add),
.data_out(VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X2n1;
wire VMR_L1D3_VMS_L1D3PHI1X2n1_wr_en;
wire [5:0] VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2_number;
wire [10:0] VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2_read_add;
wire [18:0] VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2;
VMStubs #("Tracklet") VMS_L1D3PHI1X2n1(
.data_in(VMR_L1D3_VMS_L1D3PHI1X2n1),
.enable(VMR_L1D3_VMS_L1D3PHI1X2n1_wr_en),
.number_out(VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2_number),
.read_add(VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2_read_add),
.data_out(VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI1X2n2;
wire VMR_L2D3_VMS_L2D3PHI1X2n2_wr_en;
wire [5:0] VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2_number;
wire [10:0] VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2_read_add;
wire [18:0] VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2;
VMStubs #("Tracklet") VMS_L2D3PHI1X2n2(
.data_in(VMR_L2D3_VMS_L2D3PHI1X2n2),
.enable(VMR_L2D3_VMS_L2D3PHI1X2n2_wr_en),
.number_out(VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2_number),
.read_add(VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2_read_add),
.data_out(VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X2n2;
wire VMR_L1D3_VMS_L1D3PHI1X2n2_wr_en;
wire [5:0] VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2_number;
wire [10:0] VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2_read_add;
wire [18:0] VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2;
VMStubs #("Tracklet") VMS_L1D3PHI1X2n2(
.data_in(VMR_L1D3_VMS_L1D3PHI1X2n2),
.enable(VMR_L1D3_VMS_L1D3PHI1X2n2_wr_en),
.number_out(VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2_number),
.read_add(VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2_read_add),
.data_out(VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X2n3;
wire VMR_L2D3_VMS_L2D3PHI2X2n3_wr_en;
wire [5:0] VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2_number;
wire [10:0] VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2_read_add;
wire [18:0] VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2;
VMStubs #("Tracklet") VMS_L2D3PHI2X2n3(
.data_in(VMR_L2D3_VMS_L2D3PHI2X2n3),
.enable(VMR_L2D3_VMS_L2D3PHI2X2n3_wr_en),
.number_out(VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2_number),
.read_add(VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2_read_add),
.data_out(VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X2n1;
wire VMR_L1D3_VMS_L1D3PHI2X2n1_wr_en;
wire [5:0] VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2_number;
wire [10:0] VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2_read_add;
wire [18:0] VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2;
VMStubs #("Tracklet") VMS_L1D3PHI2X2n1(
.data_in(VMR_L1D3_VMS_L1D3PHI2X2n1),
.enable(VMR_L1D3_VMS_L1D3PHI2X2n1_wr_en),
.number_out(VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2_number),
.read_add(VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2_read_add),
.data_out(VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X2n4;
wire VMR_L2D3_VMS_L2D3PHI2X2n4_wr_en;
wire [5:0] VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2_number;
wire [10:0] VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2_read_add;
wire [18:0] VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2;
VMStubs #("Tracklet") VMS_L2D3PHI2X2n4(
.data_in(VMR_L2D3_VMS_L2D3PHI2X2n4),
.enable(VMR_L2D3_VMS_L2D3PHI2X2n4_wr_en),
.number_out(VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2_number),
.read_add(VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2_read_add),
.data_out(VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X2n2;
wire VMR_L1D3_VMS_L1D3PHI2X2n2_wr_en;
wire [5:0] VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2_number;
wire [10:0] VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2_read_add;
wire [18:0] VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2;
VMStubs #("Tracklet") VMS_L1D3PHI2X2n2(
.data_in(VMR_L1D3_VMS_L1D3PHI2X2n2),
.enable(VMR_L1D3_VMS_L1D3PHI2X2n2_wr_en),
.number_out(VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2_number),
.read_add(VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2_read_add),
.data_out(VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X2n3;
wire VMR_L2D3_VMS_L2D3PHI3X2n3_wr_en;
wire [5:0] VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2_number;
wire [10:0] VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2_read_add;
wire [18:0] VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2;
VMStubs #("Tracklet") VMS_L2D3PHI3X2n3(
.data_in(VMR_L2D3_VMS_L2D3PHI3X2n3),
.enable(VMR_L2D3_VMS_L2D3PHI3X2n3_wr_en),
.number_out(VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2_number),
.read_add(VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2_read_add),
.data_out(VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X2n1;
wire VMR_L1D3_VMS_L1D3PHI3X2n1_wr_en;
wire [5:0] VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2_number;
wire [10:0] VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2_read_add;
wire [18:0] VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2;
VMStubs #("Tracklet") VMS_L1D3PHI3X2n1(
.data_in(VMR_L1D3_VMS_L1D3PHI3X2n1),
.enable(VMR_L1D3_VMS_L1D3PHI3X2n1_wr_en),
.number_out(VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2_number),
.read_add(VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2_read_add),
.data_out(VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X2n4;
wire VMR_L2D3_VMS_L2D3PHI3X2n4_wr_en;
wire [5:0] VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2_number;
wire [10:0] VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2_read_add;
wire [18:0] VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2;
VMStubs #("Tracklet") VMS_L2D3PHI3X2n4(
.data_in(VMR_L2D3_VMS_L2D3PHI3X2n4),
.enable(VMR_L2D3_VMS_L2D3PHI3X2n4_wr_en),
.number_out(VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2_number),
.read_add(VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2_read_add),
.data_out(VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X2n2;
wire VMR_L1D3_VMS_L1D3PHI3X2n2_wr_en;
wire [5:0] VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_number;
wire [10:0] VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_read_add;
wire [18:0] VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2;
VMStubs #("Tracklet") VMS_L1D3PHI3X2n2(
.data_in(VMR_L1D3_VMS_L1D3PHI3X2n2),
.enable(VMR_L1D3_VMS_L1D3PHI3X2n2_wr_en),
.number_out(VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_number),
.read_add(VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_read_add),
.data_out(VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI4X2n2;
wire VMR_L2D3_VMS_L2D3PHI4X2n2_wr_en;
wire [5:0] VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_number;
wire [10:0] VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_read_add;
wire [18:0] VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2;
VMStubs #("Tracklet") VMS_L2D3PHI4X2n2(
.data_in(VMR_L2D3_VMS_L2D3PHI4X2n2),
.enable(VMR_L2D3_VMS_L2D3PHI4X2n2_wr_en),
.number_out(VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_number),
.read_add(VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_read_add),
.data_out(VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X1n5;
wire VMR_L1D3_VMS_L1D3PHI1X1n5_wr_en;
wire [5:0] VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1_number;
wire [10:0] VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1_read_add;
wire [18:0] VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1;
VMStubs #("Tracklet") VMS_L1D3PHI1X1n5(
.data_in(VMR_L1D3_VMS_L1D3PHI1X1n5),
.enable(VMR_L1D3_VMS_L1D3PHI1X1n5_wr_en),
.number_out(VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1_number),
.read_add(VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1_read_add),
.data_out(VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI1X1n1;
wire VMR_L2D4_VMS_L2D4PHI1X1n1_wr_en;
wire [5:0] VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1_number;
wire [10:0] VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1_read_add;
wire [18:0] VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1;
VMStubs #("Tracklet") VMS_L2D4PHI1X1n1(
.data_in(VMR_L2D4_VMS_L2D4PHI1X1n1),
.enable(VMR_L2D4_VMS_L2D4PHI1X1n1_wr_en),
.number_out(VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1_number),
.read_add(VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1_read_add),
.data_out(VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X1n6;
wire VMR_L1D3_VMS_L1D3PHI1X1n6_wr_en;
wire [5:0] VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1_number;
wire [10:0] VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1_read_add;
wire [18:0] VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1;
VMStubs #("Tracklet") VMS_L1D3PHI1X1n6(
.data_in(VMR_L1D3_VMS_L1D3PHI1X1n6),
.enable(VMR_L1D3_VMS_L1D3PHI1X1n6_wr_en),
.number_out(VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1_number),
.read_add(VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1_read_add),
.data_out(VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X1n1;
wire VMR_L2D4_VMS_L2D4PHI2X1n1_wr_en;
wire [5:0] VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1_number;
wire [10:0] VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1_read_add;
wire [18:0] VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1;
VMStubs #("Tracklet") VMS_L2D4PHI2X1n1(
.data_in(VMR_L2D4_VMS_L2D4PHI2X1n1),
.enable(VMR_L2D4_VMS_L2D4PHI2X1n1_wr_en),
.number_out(VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1_number),
.read_add(VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1_read_add),
.data_out(VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X1n5;
wire VMR_L1D3_VMS_L1D3PHI2X1n5_wr_en;
wire [5:0] VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1_number;
wire [10:0] VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1_read_add;
wire [18:0] VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1;
VMStubs #("Tracklet") VMS_L1D3PHI2X1n5(
.data_in(VMR_L1D3_VMS_L1D3PHI2X1n5),
.enable(VMR_L1D3_VMS_L1D3PHI2X1n5_wr_en),
.number_out(VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1_number),
.read_add(VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1_read_add),
.data_out(VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X1n2;
wire VMR_L2D4_VMS_L2D4PHI2X1n2_wr_en;
wire [5:0] VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1_number;
wire [10:0] VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1_read_add;
wire [18:0] VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1;
VMStubs #("Tracklet") VMS_L2D4PHI2X1n2(
.data_in(VMR_L2D4_VMS_L2D4PHI2X1n2),
.enable(VMR_L2D4_VMS_L2D4PHI2X1n2_wr_en),
.number_out(VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1_number),
.read_add(VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1_read_add),
.data_out(VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X1n6;
wire VMR_L1D3_VMS_L1D3PHI2X1n6_wr_en;
wire [5:0] VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1_number;
wire [10:0] VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1_read_add;
wire [18:0] VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1;
VMStubs #("Tracklet") VMS_L1D3PHI2X1n6(
.data_in(VMR_L1D3_VMS_L1D3PHI2X1n6),
.enable(VMR_L1D3_VMS_L1D3PHI2X1n6_wr_en),
.number_out(VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1_number),
.read_add(VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1_read_add),
.data_out(VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X1n1;
wire VMR_L2D4_VMS_L2D4PHI3X1n1_wr_en;
wire [5:0] VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1_number;
wire [10:0] VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1_read_add;
wire [18:0] VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1;
VMStubs #("Tracklet") VMS_L2D4PHI3X1n1(
.data_in(VMR_L2D4_VMS_L2D4PHI3X1n1),
.enable(VMR_L2D4_VMS_L2D4PHI3X1n1_wr_en),
.number_out(VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1_number),
.read_add(VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1_read_add),
.data_out(VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X1n5;
wire VMR_L1D3_VMS_L1D3PHI3X1n5_wr_en;
wire [5:0] VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1_number;
wire [10:0] VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1_read_add;
wire [18:0] VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1;
VMStubs #("Tracklet") VMS_L1D3PHI3X1n5(
.data_in(VMR_L1D3_VMS_L1D3PHI3X1n5),
.enable(VMR_L1D3_VMS_L1D3PHI3X1n5_wr_en),
.number_out(VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1_number),
.read_add(VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1_read_add),
.data_out(VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X1n2;
wire VMR_L2D4_VMS_L2D4PHI3X1n2_wr_en;
wire [5:0] VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1_number;
wire [10:0] VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1_read_add;
wire [18:0] VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1;
VMStubs #("Tracklet") VMS_L2D4PHI3X1n2(
.data_in(VMR_L2D4_VMS_L2D4PHI3X1n2),
.enable(VMR_L2D4_VMS_L2D4PHI3X1n2_wr_en),
.number_out(VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1_number),
.read_add(VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1_read_add),
.data_out(VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X1n6;
wire VMR_L1D3_VMS_L1D3PHI3X1n6_wr_en;
wire [5:0] VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1_number;
wire [10:0] VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1_read_add;
wire [18:0] VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1;
VMStubs #("Tracklet") VMS_L1D3PHI3X1n6(
.data_in(VMR_L1D3_VMS_L1D3PHI3X1n6),
.enable(VMR_L1D3_VMS_L1D3PHI3X1n6_wr_en),
.number_out(VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1_number),
.read_add(VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1_read_add),
.data_out(VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI4X1n1;
wire VMR_L2D4_VMS_L2D4PHI4X1n1_wr_en;
wire [5:0] VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1_number;
wire [10:0] VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1_read_add;
wire [18:0] VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1;
VMStubs #("Tracklet") VMS_L2D4PHI4X1n1(
.data_in(VMR_L2D4_VMS_L2D4PHI4X1n1),
.enable(VMR_L2D4_VMS_L2D4PHI4X1n1_wr_en),
.number_out(VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1_number),
.read_add(VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1_read_add),
.data_out(VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X2n3;
wire VMR_L1D3_VMS_L1D3PHI1X2n3_wr_en;
wire [5:0] VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1_number;
wire [10:0] VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1_read_add;
wire [18:0] VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1;
VMStubs #("Tracklet") VMS_L1D3PHI1X2n3(
.data_in(VMR_L1D3_VMS_L1D3PHI1X2n3),
.enable(VMR_L1D3_VMS_L1D3PHI1X2n3_wr_en),
.number_out(VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1_number),
.read_add(VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1_read_add),
.data_out(VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI1X1n2;
wire VMR_L2D4_VMS_L2D4PHI1X1n2_wr_en;
wire [5:0] VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1_number;
wire [10:0] VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1_read_add;
wire [18:0] VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1;
VMStubs #("Tracklet") VMS_L2D4PHI1X1n2(
.data_in(VMR_L2D4_VMS_L2D4PHI1X1n2),
.enable(VMR_L2D4_VMS_L2D4PHI1X1n2_wr_en),
.number_out(VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1_number),
.read_add(VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1_read_add),
.data_out(VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X2n4;
wire VMR_L1D3_VMS_L1D3PHI1X2n4_wr_en;
wire [5:0] VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1_number;
wire [10:0] VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1_read_add;
wire [18:0] VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1;
VMStubs #("Tracklet") VMS_L1D3PHI1X2n4(
.data_in(VMR_L1D3_VMS_L1D3PHI1X2n4),
.enable(VMR_L1D3_VMS_L1D3PHI1X2n4_wr_en),
.number_out(VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1_number),
.read_add(VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1_read_add),
.data_out(VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X1n3;
wire VMR_L2D4_VMS_L2D4PHI2X1n3_wr_en;
wire [5:0] VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1_number;
wire [10:0] VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1_read_add;
wire [18:0] VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1;
VMStubs #("Tracklet") VMS_L2D4PHI2X1n3(
.data_in(VMR_L2D4_VMS_L2D4PHI2X1n3),
.enable(VMR_L2D4_VMS_L2D4PHI2X1n3_wr_en),
.number_out(VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1_number),
.read_add(VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1_read_add),
.data_out(VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X2n3;
wire VMR_L1D3_VMS_L1D3PHI2X2n3_wr_en;
wire [5:0] VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1_number;
wire [10:0] VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1_read_add;
wire [18:0] VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1;
VMStubs #("Tracklet") VMS_L1D3PHI2X2n3(
.data_in(VMR_L1D3_VMS_L1D3PHI2X2n3),
.enable(VMR_L1D3_VMS_L1D3PHI2X2n3_wr_en),
.number_out(VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1_number),
.read_add(VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1_read_add),
.data_out(VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X1n4;
wire VMR_L2D4_VMS_L2D4PHI2X1n4_wr_en;
wire [5:0] VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1_number;
wire [10:0] VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1_read_add;
wire [18:0] VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1;
VMStubs #("Tracklet") VMS_L2D4PHI2X1n4(
.data_in(VMR_L2D4_VMS_L2D4PHI2X1n4),
.enable(VMR_L2D4_VMS_L2D4PHI2X1n4_wr_en),
.number_out(VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1_number),
.read_add(VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1_read_add),
.data_out(VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X2n4;
wire VMR_L1D3_VMS_L1D3PHI2X2n4_wr_en;
wire [5:0] VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1_number;
wire [10:0] VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1_read_add;
wire [18:0] VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1;
VMStubs #("Tracklet") VMS_L1D3PHI2X2n4(
.data_in(VMR_L1D3_VMS_L1D3PHI2X2n4),
.enable(VMR_L1D3_VMS_L1D3PHI2X2n4_wr_en),
.number_out(VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1_number),
.read_add(VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1_read_add),
.data_out(VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X1n3;
wire VMR_L2D4_VMS_L2D4PHI3X1n3_wr_en;
wire [5:0] VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1_number;
wire [10:0] VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1_read_add;
wire [18:0] VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1;
VMStubs #("Tracklet") VMS_L2D4PHI3X1n3(
.data_in(VMR_L2D4_VMS_L2D4PHI3X1n3),
.enable(VMR_L2D4_VMS_L2D4PHI3X1n3_wr_en),
.number_out(VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1_number),
.read_add(VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1_read_add),
.data_out(VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X2n3;
wire VMR_L1D3_VMS_L1D3PHI3X2n3_wr_en;
wire [5:0] VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1_number;
wire [10:0] VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1_read_add;
wire [18:0] VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1;
VMStubs #("Tracklet") VMS_L1D3PHI3X2n3(
.data_in(VMR_L1D3_VMS_L1D3PHI3X2n3),
.enable(VMR_L1D3_VMS_L1D3PHI3X2n3_wr_en),
.number_out(VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1_number),
.read_add(VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1_read_add),
.data_out(VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X1n4;
wire VMR_L2D4_VMS_L2D4PHI3X1n4_wr_en;
wire [5:0] VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1_number;
wire [10:0] VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1_read_add;
wire [18:0] VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1;
VMStubs #("Tracklet") VMS_L2D4PHI3X1n4(
.data_in(VMR_L2D4_VMS_L2D4PHI3X1n4),
.enable(VMR_L2D4_VMS_L2D4PHI3X1n4_wr_en),
.number_out(VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1_number),
.read_add(VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1_read_add),
.data_out(VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X2n4;
wire VMR_L1D3_VMS_L1D3PHI3X2n4_wr_en;
wire [5:0] VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1_number;
wire [10:0] VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1_read_add;
wire [18:0] VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1;
VMStubs #("Tracklet") VMS_L1D3PHI3X2n4(
.data_in(VMR_L1D3_VMS_L1D3PHI3X2n4),
.enable(VMR_L1D3_VMS_L1D3PHI3X2n4_wr_en),
.number_out(VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1_number),
.read_add(VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1_read_add),
.data_out(VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI4X1n2;
wire VMR_L2D4_VMS_L2D4PHI4X1n2_wr_en;
wire [5:0] VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1_number;
wire [10:0] VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1_read_add;
wire [18:0] VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1;
VMStubs #("Tracklet") VMS_L2D4PHI4X1n2(
.data_in(VMR_L2D4_VMS_L2D4PHI4X1n2),
.enable(VMR_L2D4_VMS_L2D4PHI4X1n2_wr_en),
.number_out(VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1_number),
.read_add(VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1_read_add),
.data_out(VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X2n5;
wire VMR_L1D3_VMS_L1D3PHI1X2n5_wr_en;
wire [5:0] VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2_number;
wire [10:0] VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2_read_add;
wire [18:0] VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2;
VMStubs #("Tracklet") VMS_L1D3PHI1X2n5(
.data_in(VMR_L1D3_VMS_L1D3PHI1X2n5),
.enable(VMR_L1D3_VMS_L1D3PHI1X2n5_wr_en),
.number_out(VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2_number),
.read_add(VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2_read_add),
.data_out(VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI1X2n1;
wire VMR_L2D4_VMS_L2D4PHI1X2n1_wr_en;
wire [5:0] VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2_number;
wire [10:0] VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2_read_add;
wire [18:0] VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2;
VMStubs #("Tracklet") VMS_L2D4PHI1X2n1(
.data_in(VMR_L2D4_VMS_L2D4PHI1X2n1),
.enable(VMR_L2D4_VMS_L2D4PHI1X2n1_wr_en),
.number_out(VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2_number),
.read_add(VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2_read_add),
.data_out(VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X2n6;
wire VMR_L1D3_VMS_L1D3PHI1X2n6_wr_en;
wire [5:0] VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2_number;
wire [10:0] VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2_read_add;
wire [18:0] VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2;
VMStubs #("Tracklet") VMS_L1D3PHI1X2n6(
.data_in(VMR_L1D3_VMS_L1D3PHI1X2n6),
.enable(VMR_L1D3_VMS_L1D3PHI1X2n6_wr_en),
.number_out(VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2_number),
.read_add(VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2_read_add),
.data_out(VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X2n1;
wire VMR_L2D4_VMS_L2D4PHI2X2n1_wr_en;
wire [5:0] VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2_number;
wire [10:0] VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2_read_add;
wire [18:0] VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2;
VMStubs #("Tracklet") VMS_L2D4PHI2X2n1(
.data_in(VMR_L2D4_VMS_L2D4PHI2X2n1),
.enable(VMR_L2D4_VMS_L2D4PHI2X2n1_wr_en),
.number_out(VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2_number),
.read_add(VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2_read_add),
.data_out(VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X2n5;
wire VMR_L1D3_VMS_L1D3PHI2X2n5_wr_en;
wire [5:0] VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2_number;
wire [10:0] VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2_read_add;
wire [18:0] VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2;
VMStubs #("Tracklet") VMS_L1D3PHI2X2n5(
.data_in(VMR_L1D3_VMS_L1D3PHI2X2n5),
.enable(VMR_L1D3_VMS_L1D3PHI2X2n5_wr_en),
.number_out(VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2_number),
.read_add(VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2_read_add),
.data_out(VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X2n2;
wire VMR_L2D4_VMS_L2D4PHI2X2n2_wr_en;
wire [5:0] VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2_number;
wire [10:0] VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2_read_add;
wire [18:0] VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2;
VMStubs #("Tracklet") VMS_L2D4PHI2X2n2(
.data_in(VMR_L2D4_VMS_L2D4PHI2X2n2),
.enable(VMR_L2D4_VMS_L2D4PHI2X2n2_wr_en),
.number_out(VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2_number),
.read_add(VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2_read_add),
.data_out(VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X2n6;
wire VMR_L1D3_VMS_L1D3PHI2X2n6_wr_en;
wire [5:0] VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2_number;
wire [10:0] VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2_read_add;
wire [18:0] VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2;
VMStubs #("Tracklet") VMS_L1D3PHI2X2n6(
.data_in(VMR_L1D3_VMS_L1D3PHI2X2n6),
.enable(VMR_L1D3_VMS_L1D3PHI2X2n6_wr_en),
.number_out(VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2_number),
.read_add(VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2_read_add),
.data_out(VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X2n1;
wire VMR_L2D4_VMS_L2D4PHI3X2n1_wr_en;
wire [5:0] VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2_number;
wire [10:0] VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2_read_add;
wire [18:0] VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2;
VMStubs #("Tracklet") VMS_L2D4PHI3X2n1(
.data_in(VMR_L2D4_VMS_L2D4PHI3X2n1),
.enable(VMR_L2D4_VMS_L2D4PHI3X2n1_wr_en),
.number_out(VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2_number),
.read_add(VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2_read_add),
.data_out(VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X2n5;
wire VMR_L1D3_VMS_L1D3PHI3X2n5_wr_en;
wire [5:0] VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2_number;
wire [10:0] VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2_read_add;
wire [18:0] VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2;
VMStubs #("Tracklet") VMS_L1D3PHI3X2n5(
.data_in(VMR_L1D3_VMS_L1D3PHI3X2n5),
.enable(VMR_L1D3_VMS_L1D3PHI3X2n5_wr_en),
.number_out(VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2_number),
.read_add(VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2_read_add),
.data_out(VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X2n2;
wire VMR_L2D4_VMS_L2D4PHI3X2n2_wr_en;
wire [5:0] VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2_number;
wire [10:0] VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2_read_add;
wire [18:0] VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2;
VMStubs #("Tracklet") VMS_L2D4PHI3X2n2(
.data_in(VMR_L2D4_VMS_L2D4PHI3X2n2),
.enable(VMR_L2D4_VMS_L2D4PHI3X2n2_wr_en),
.number_out(VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2_number),
.read_add(VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2_read_add),
.data_out(VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X2n6;
wire VMR_L1D3_VMS_L1D3PHI3X2n6_wr_en;
wire [5:0] VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2_number;
wire [10:0] VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2_read_add;
wire [18:0] VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2;
VMStubs #("Tracklet") VMS_L1D3PHI3X2n6(
.data_in(VMR_L1D3_VMS_L1D3PHI3X2n6),
.enable(VMR_L1D3_VMS_L1D3PHI3X2n6_wr_en),
.number_out(VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2_number),
.read_add(VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2_read_add),
.data_out(VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI4X2n1;
wire VMR_L2D4_VMS_L2D4PHI4X2n1_wr_en;
wire [5:0] VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2_number;
wire [10:0] VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2_read_add;
wire [18:0] VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2;
VMStubs #("Tracklet") VMS_L2D4PHI4X2n1(
.data_in(VMR_L2D4_VMS_L2D4PHI4X2n1),
.enable(VMR_L2D4_VMS_L2D4PHI4X2n1_wr_en),
.number_out(VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2_number),
.read_add(VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2_read_add),
.data_out(VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI1X1n1;
wire VMR_L1D4_VMS_L1D4PHI1X1n1_wr_en;
wire [5:0] VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2_number;
wire [10:0] VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2_read_add;
wire [18:0] VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2;
VMStubs #("Tracklet") VMS_L1D4PHI1X1n1(
.data_in(VMR_L1D4_VMS_L1D4PHI1X1n1),
.enable(VMR_L1D4_VMS_L1D4PHI1X1n1_wr_en),
.number_out(VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2_number),
.read_add(VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2_read_add),
.data_out(VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI1X2n2;
wire VMR_L2D4_VMS_L2D4PHI1X2n2_wr_en;
wire [5:0] VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2_number;
wire [10:0] VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2_read_add;
wire [18:0] VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2;
VMStubs #("Tracklet") VMS_L2D4PHI1X2n2(
.data_in(VMR_L2D4_VMS_L2D4PHI1X2n2),
.enable(VMR_L2D4_VMS_L2D4PHI1X2n2_wr_en),
.number_out(VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2_number),
.read_add(VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2_read_add),
.data_out(VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI1X1n2;
wire VMR_L1D4_VMS_L1D4PHI1X1n2_wr_en;
wire [5:0] VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2_number;
wire [10:0] VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2_read_add;
wire [18:0] VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2;
VMStubs #("Tracklet") VMS_L1D4PHI1X1n2(
.data_in(VMR_L1D4_VMS_L1D4PHI1X1n2),
.enable(VMR_L1D4_VMS_L1D4PHI1X1n2_wr_en),
.number_out(VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2_number),
.read_add(VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2_read_add),
.data_out(VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X2n3;
wire VMR_L2D4_VMS_L2D4PHI2X2n3_wr_en;
wire [5:0] VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2_number;
wire [10:0] VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2_read_add;
wire [18:0] VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2;
VMStubs #("Tracklet") VMS_L2D4PHI2X2n3(
.data_in(VMR_L2D4_VMS_L2D4PHI2X2n3),
.enable(VMR_L2D4_VMS_L2D4PHI2X2n3_wr_en),
.number_out(VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2_number),
.read_add(VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2_read_add),
.data_out(VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI2X1n1;
wire VMR_L1D4_VMS_L1D4PHI2X1n1_wr_en;
wire [5:0] VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2_number;
wire [10:0] VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2_read_add;
wire [18:0] VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2;
VMStubs #("Tracklet") VMS_L1D4PHI2X1n1(
.data_in(VMR_L1D4_VMS_L1D4PHI2X1n1),
.enable(VMR_L1D4_VMS_L1D4PHI2X1n1_wr_en),
.number_out(VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2_number),
.read_add(VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2_read_add),
.data_out(VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X2n4;
wire VMR_L2D4_VMS_L2D4PHI2X2n4_wr_en;
wire [5:0] VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2_number;
wire [10:0] VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2_read_add;
wire [18:0] VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2;
VMStubs #("Tracklet") VMS_L2D4PHI2X2n4(
.data_in(VMR_L2D4_VMS_L2D4PHI2X2n4),
.enable(VMR_L2D4_VMS_L2D4PHI2X2n4_wr_en),
.number_out(VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2_number),
.read_add(VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2_read_add),
.data_out(VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI2X1n2;
wire VMR_L1D4_VMS_L1D4PHI2X1n2_wr_en;
wire [5:0] VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2_number;
wire [10:0] VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2_read_add;
wire [18:0] VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2;
VMStubs #("Tracklet") VMS_L1D4PHI2X1n2(
.data_in(VMR_L1D4_VMS_L1D4PHI2X1n2),
.enable(VMR_L1D4_VMS_L1D4PHI2X1n2_wr_en),
.number_out(VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2_number),
.read_add(VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2_read_add),
.data_out(VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X2n3;
wire VMR_L2D4_VMS_L2D4PHI3X2n3_wr_en;
wire [5:0] VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2_number;
wire [10:0] VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2_read_add;
wire [18:0] VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2;
VMStubs #("Tracklet") VMS_L2D4PHI3X2n3(
.data_in(VMR_L2D4_VMS_L2D4PHI3X2n3),
.enable(VMR_L2D4_VMS_L2D4PHI3X2n3_wr_en),
.number_out(VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2_number),
.read_add(VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2_read_add),
.data_out(VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI3X1n1;
wire VMR_L1D4_VMS_L1D4PHI3X1n1_wr_en;
wire [5:0] VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2_number;
wire [10:0] VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2_read_add;
wire [18:0] VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2;
VMStubs #("Tracklet") VMS_L1D4PHI3X1n1(
.data_in(VMR_L1D4_VMS_L1D4PHI3X1n1),
.enable(VMR_L1D4_VMS_L1D4PHI3X1n1_wr_en),
.number_out(VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2_number),
.read_add(VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2_read_add),
.data_out(VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X2n4;
wire VMR_L2D4_VMS_L2D4PHI3X2n4_wr_en;
wire [5:0] VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2_number;
wire [10:0] VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2_read_add;
wire [18:0] VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2;
VMStubs #("Tracklet") VMS_L2D4PHI3X2n4(
.data_in(VMR_L2D4_VMS_L2D4PHI3X2n4),
.enable(VMR_L2D4_VMS_L2D4PHI3X2n4_wr_en),
.number_out(VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2_number),
.read_add(VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2_read_add),
.data_out(VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI3X1n2;
wire VMR_L1D4_VMS_L1D4PHI3X1n2_wr_en;
wire [5:0] VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2_number;
wire [10:0] VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2_read_add;
wire [18:0] VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2;
VMStubs #("Tracklet") VMS_L1D4PHI3X1n2(
.data_in(VMR_L1D4_VMS_L1D4PHI3X1n2),
.enable(VMR_L1D4_VMS_L1D4PHI3X1n2_wr_en),
.number_out(VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2_number),
.read_add(VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2_read_add),
.data_out(VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI4X2n2;
wire VMR_L2D4_VMS_L2D4PHI4X2n2_wr_en;
wire [5:0] VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2_number;
wire [10:0] VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2_read_add;
wire [18:0] VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2;
VMStubs #("Tracklet") VMS_L2D4PHI4X2n2(
.data_in(VMR_L2D4_VMS_L2D4PHI4X2n2),
.enable(VMR_L2D4_VMS_L2D4PHI4X2n2_wr_en),
.number_out(VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2_number),
.read_add(VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2_read_add),
.data_out(VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X1n1;
wire VMR_L3D3_VMS_L3D3PHI1X1n1_wr_en;
wire [5:0] VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_number;
wire [10:0] VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_read_add;
wire [18:0] VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1;
VMStubs #("Tracklet") VMS_L3D3PHI1X1n1(
.data_in(VMR_L3D3_VMS_L3D3PHI1X1n1),
.enable(VMR_L3D3_VMS_L3D3PHI1X1n1_wr_en),
.number_out(VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_number),
.read_add(VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_read_add),
.data_out(VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI1X1n1;
wire VMR_L4D3_VMS_L4D3PHI1X1n1_wr_en;
wire [5:0] VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_number;
wire [10:0] VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_read_add;
wire [18:0] VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1;
VMStubs #("Tracklet") VMS_L4D3PHI1X1n1(
.data_in(VMR_L4D3_VMS_L4D3PHI1X1n1),
.enable(VMR_L4D3_VMS_L4D3PHI1X1n1_wr_en),
.number_out(VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_number),
.read_add(VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_read_add),
.data_out(VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X1n2;
wire VMR_L3D3_VMS_L3D3PHI1X1n2_wr_en;
wire [5:0] VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1_number;
wire [10:0] VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1_read_add;
wire [18:0] VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1;
VMStubs #("Tracklet") VMS_L3D3PHI1X1n2(
.data_in(VMR_L3D3_VMS_L3D3PHI1X1n2),
.enable(VMR_L3D3_VMS_L3D3PHI1X1n2_wr_en),
.number_out(VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1_number),
.read_add(VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1_read_add),
.data_out(VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X1n1;
wire VMR_L4D3_VMS_L4D3PHI2X1n1_wr_en;
wire [5:0] VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1_number;
wire [10:0] VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1_read_add;
wire [18:0] VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1;
VMStubs #("Tracklet") VMS_L4D3PHI2X1n1(
.data_in(VMR_L4D3_VMS_L4D3PHI2X1n1),
.enable(VMR_L4D3_VMS_L4D3PHI2X1n1_wr_en),
.number_out(VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1_number),
.read_add(VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1_read_add),
.data_out(VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X1n1;
wire VMR_L3D3_VMS_L3D3PHI2X1n1_wr_en;
wire [5:0] VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1_number;
wire [10:0] VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1_read_add;
wire [18:0] VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1;
VMStubs #("Tracklet") VMS_L3D3PHI2X1n1(
.data_in(VMR_L3D3_VMS_L3D3PHI2X1n1),
.enable(VMR_L3D3_VMS_L3D3PHI2X1n1_wr_en),
.number_out(VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1_number),
.read_add(VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1_read_add),
.data_out(VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X1n2;
wire VMR_L4D3_VMS_L4D3PHI2X1n2_wr_en;
wire [5:0] VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1_number;
wire [10:0] VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1_read_add;
wire [18:0] VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1;
VMStubs #("Tracklet") VMS_L4D3PHI2X1n2(
.data_in(VMR_L4D3_VMS_L4D3PHI2X1n2),
.enable(VMR_L4D3_VMS_L4D3PHI2X1n2_wr_en),
.number_out(VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1_number),
.read_add(VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1_read_add),
.data_out(VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X1n2;
wire VMR_L3D3_VMS_L3D3PHI2X1n2_wr_en;
wire [5:0] VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1_number;
wire [10:0] VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1_read_add;
wire [18:0] VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1;
VMStubs #("Tracklet") VMS_L3D3PHI2X1n2(
.data_in(VMR_L3D3_VMS_L3D3PHI2X1n2),
.enable(VMR_L3D3_VMS_L3D3PHI2X1n2_wr_en),
.number_out(VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1_number),
.read_add(VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1_read_add),
.data_out(VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X1n1;
wire VMR_L4D3_VMS_L4D3PHI3X1n1_wr_en;
wire [5:0] VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1_number;
wire [10:0] VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1_read_add;
wire [18:0] VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1;
VMStubs #("Tracklet") VMS_L4D3PHI3X1n1(
.data_in(VMR_L4D3_VMS_L4D3PHI3X1n1),
.enable(VMR_L4D3_VMS_L4D3PHI3X1n1_wr_en),
.number_out(VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1_number),
.read_add(VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1_read_add),
.data_out(VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X1n1;
wire VMR_L3D3_VMS_L3D3PHI3X1n1_wr_en;
wire [5:0] VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1_number;
wire [10:0] VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1_read_add;
wire [18:0] VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1;
VMStubs #("Tracklet") VMS_L3D3PHI3X1n1(
.data_in(VMR_L3D3_VMS_L3D3PHI3X1n1),
.enable(VMR_L3D3_VMS_L3D3PHI3X1n1_wr_en),
.number_out(VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1_number),
.read_add(VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1_read_add),
.data_out(VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X1n2;
wire VMR_L4D3_VMS_L4D3PHI3X1n2_wr_en;
wire [5:0] VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1_number;
wire [10:0] VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1_read_add;
wire [18:0] VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1;
VMStubs #("Tracklet") VMS_L4D3PHI3X1n2(
.data_in(VMR_L4D3_VMS_L4D3PHI3X1n2),
.enable(VMR_L4D3_VMS_L4D3PHI3X1n2_wr_en),
.number_out(VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1_number),
.read_add(VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1_read_add),
.data_out(VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X1n2;
wire VMR_L3D3_VMS_L3D3PHI3X1n2_wr_en;
wire [5:0] VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1_number;
wire [10:0] VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1_read_add;
wire [18:0] VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1;
VMStubs #("Tracklet") VMS_L3D3PHI3X1n2(
.data_in(VMR_L3D3_VMS_L3D3PHI3X1n2),
.enable(VMR_L3D3_VMS_L3D3PHI3X1n2_wr_en),
.number_out(VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1_number),
.read_add(VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1_read_add),
.data_out(VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI4X1n1;
wire VMR_L4D3_VMS_L4D3PHI4X1n1_wr_en;
wire [5:0] VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1_number;
wire [10:0] VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1_read_add;
wire [18:0] VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1;
VMStubs #("Tracklet") VMS_L4D3PHI4X1n1(
.data_in(VMR_L4D3_VMS_L4D3PHI4X1n1),
.enable(VMR_L4D3_VMS_L4D3PHI4X1n1_wr_en),
.number_out(VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1_number),
.read_add(VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1_read_add),
.data_out(VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X2n1;
wire VMR_L3D3_VMS_L3D3PHI1X2n1_wr_en;
wire [5:0] VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_number;
wire [10:0] VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_read_add;
wire [18:0] VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2;
VMStubs #("Tracklet") VMS_L3D3PHI1X2n1(
.data_in(VMR_L3D3_VMS_L3D3PHI1X2n1),
.enable(VMR_L3D3_VMS_L3D3PHI1X2n1_wr_en),
.number_out(VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_number),
.read_add(VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_read_add),
.data_out(VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI1X2n1;
wire VMR_L4D3_VMS_L4D3PHI1X2n1_wr_en;
wire [5:0] VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_number;
wire [10:0] VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_read_add;
wire [18:0] VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2;
VMStubs #("Tracklet") VMS_L4D3PHI1X2n1(
.data_in(VMR_L4D3_VMS_L4D3PHI1X2n1),
.enable(VMR_L4D3_VMS_L4D3PHI1X2n1_wr_en),
.number_out(VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_number),
.read_add(VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_read_add),
.data_out(VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X2n2;
wire VMR_L3D3_VMS_L3D3PHI1X2n2_wr_en;
wire [5:0] VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2_number;
wire [10:0] VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2_read_add;
wire [18:0] VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2;
VMStubs #("Tracklet") VMS_L3D3PHI1X2n2(
.data_in(VMR_L3D3_VMS_L3D3PHI1X2n2),
.enable(VMR_L3D3_VMS_L3D3PHI1X2n2_wr_en),
.number_out(VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2_number),
.read_add(VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2_read_add),
.data_out(VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X2n1;
wire VMR_L4D3_VMS_L4D3PHI2X2n1_wr_en;
wire [5:0] VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2_number;
wire [10:0] VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2_read_add;
wire [18:0] VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2;
VMStubs #("Tracklet") VMS_L4D3PHI2X2n1(
.data_in(VMR_L4D3_VMS_L4D3PHI2X2n1),
.enable(VMR_L4D3_VMS_L4D3PHI2X2n1_wr_en),
.number_out(VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2_number),
.read_add(VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2_read_add),
.data_out(VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X2n1;
wire VMR_L3D3_VMS_L3D3PHI2X2n1_wr_en;
wire [5:0] VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2_number;
wire [10:0] VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2_read_add;
wire [18:0] VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2;
VMStubs #("Tracklet") VMS_L3D3PHI2X2n1(
.data_in(VMR_L3D3_VMS_L3D3PHI2X2n1),
.enable(VMR_L3D3_VMS_L3D3PHI2X2n1_wr_en),
.number_out(VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2_number),
.read_add(VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2_read_add),
.data_out(VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X2n2;
wire VMR_L4D3_VMS_L4D3PHI2X2n2_wr_en;
wire [5:0] VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2_number;
wire [10:0] VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2_read_add;
wire [18:0] VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2;
VMStubs #("Tracklet") VMS_L4D3PHI2X2n2(
.data_in(VMR_L4D3_VMS_L4D3PHI2X2n2),
.enable(VMR_L4D3_VMS_L4D3PHI2X2n2_wr_en),
.number_out(VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2_number),
.read_add(VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2_read_add),
.data_out(VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X2n2;
wire VMR_L3D3_VMS_L3D3PHI2X2n2_wr_en;
wire [5:0] VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2_number;
wire [10:0] VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2_read_add;
wire [18:0] VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2;
VMStubs #("Tracklet") VMS_L3D3PHI2X2n2(
.data_in(VMR_L3D3_VMS_L3D3PHI2X2n2),
.enable(VMR_L3D3_VMS_L3D3PHI2X2n2_wr_en),
.number_out(VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2_number),
.read_add(VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2_read_add),
.data_out(VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X2n1;
wire VMR_L4D3_VMS_L4D3PHI3X2n1_wr_en;
wire [5:0] VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2_number;
wire [10:0] VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2_read_add;
wire [18:0] VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2;
VMStubs #("Tracklet") VMS_L4D3PHI3X2n1(
.data_in(VMR_L4D3_VMS_L4D3PHI3X2n1),
.enable(VMR_L4D3_VMS_L4D3PHI3X2n1_wr_en),
.number_out(VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2_number),
.read_add(VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2_read_add),
.data_out(VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X2n1;
wire VMR_L3D3_VMS_L3D3PHI3X2n1_wr_en;
wire [5:0] VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2_number;
wire [10:0] VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2_read_add;
wire [18:0] VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2;
VMStubs #("Tracklet") VMS_L3D3PHI3X2n1(
.data_in(VMR_L3D3_VMS_L3D3PHI3X2n1),
.enable(VMR_L3D3_VMS_L3D3PHI3X2n1_wr_en),
.number_out(VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2_number),
.read_add(VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2_read_add),
.data_out(VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X2n2;
wire VMR_L4D3_VMS_L4D3PHI3X2n2_wr_en;
wire [5:0] VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2_number;
wire [10:0] VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2_read_add;
wire [18:0] VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2;
VMStubs #("Tracklet") VMS_L4D3PHI3X2n2(
.data_in(VMR_L4D3_VMS_L4D3PHI3X2n2),
.enable(VMR_L4D3_VMS_L4D3PHI3X2n2_wr_en),
.number_out(VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2_number),
.read_add(VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2_read_add),
.data_out(VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X2n2;
wire VMR_L3D3_VMS_L3D3PHI3X2n2_wr_en;
wire [5:0] VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2_number;
wire [10:0] VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2_read_add;
wire [18:0] VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2;
VMStubs #("Tracklet") VMS_L3D3PHI3X2n2(
.data_in(VMR_L3D3_VMS_L3D3PHI3X2n2),
.enable(VMR_L3D3_VMS_L3D3PHI3X2n2_wr_en),
.number_out(VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2_number),
.read_add(VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2_read_add),
.data_out(VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI4X2n1;
wire VMR_L4D3_VMS_L4D3PHI4X2n1_wr_en;
wire [5:0] VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2_number;
wire [10:0] VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2_read_add;
wire [18:0] VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2;
VMStubs #("Tracklet") VMS_L4D3PHI4X2n1(
.data_in(VMR_L4D3_VMS_L4D3PHI4X2n1),
.enable(VMR_L4D3_VMS_L4D3PHI4X2n1_wr_en),
.number_out(VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2_number),
.read_add(VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2_read_add),
.data_out(VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X1n3;
wire VMR_L3D3_VMS_L3D3PHI1X1n3_wr_en;
wire [5:0] VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2_number;
wire [10:0] VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2_read_add;
wire [18:0] VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2;
VMStubs #("Tracklet") VMS_L3D3PHI1X1n3(
.data_in(VMR_L3D3_VMS_L3D3PHI1X1n3),
.enable(VMR_L3D3_VMS_L3D3PHI1X1n3_wr_en),
.number_out(VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2_number),
.read_add(VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2_read_add),
.data_out(VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI1X2n2;
wire VMR_L4D3_VMS_L4D3PHI1X2n2_wr_en;
wire [5:0] VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2_number;
wire [10:0] VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2_read_add;
wire [18:0] VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2;
VMStubs #("Tracklet") VMS_L4D3PHI1X2n2(
.data_in(VMR_L4D3_VMS_L4D3PHI1X2n2),
.enable(VMR_L4D3_VMS_L4D3PHI1X2n2_wr_en),
.number_out(VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2_number),
.read_add(VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2_read_add),
.data_out(VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X1n4;
wire VMR_L3D3_VMS_L3D3PHI1X1n4_wr_en;
wire [5:0] VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2_number;
wire [10:0] VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2_read_add;
wire [18:0] VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2;
VMStubs #("Tracklet") VMS_L3D3PHI1X1n4(
.data_in(VMR_L3D3_VMS_L3D3PHI1X1n4),
.enable(VMR_L3D3_VMS_L3D3PHI1X1n4_wr_en),
.number_out(VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2_number),
.read_add(VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2_read_add),
.data_out(VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X2n3;
wire VMR_L4D3_VMS_L4D3PHI2X2n3_wr_en;
wire [5:0] VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2_number;
wire [10:0] VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2_read_add;
wire [18:0] VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2;
VMStubs #("Tracklet") VMS_L4D3PHI2X2n3(
.data_in(VMR_L4D3_VMS_L4D3PHI2X2n3),
.enable(VMR_L4D3_VMS_L4D3PHI2X2n3_wr_en),
.number_out(VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2_number),
.read_add(VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2_read_add),
.data_out(VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X1n3;
wire VMR_L3D3_VMS_L3D3PHI2X1n3_wr_en;
wire [5:0] VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2_number;
wire [10:0] VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2_read_add;
wire [18:0] VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2;
VMStubs #("Tracklet") VMS_L3D3PHI2X1n3(
.data_in(VMR_L3D3_VMS_L3D3PHI2X1n3),
.enable(VMR_L3D3_VMS_L3D3PHI2X1n3_wr_en),
.number_out(VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2_number),
.read_add(VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2_read_add),
.data_out(VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X2n4;
wire VMR_L4D3_VMS_L4D3PHI2X2n4_wr_en;
wire [5:0] VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2_number;
wire [10:0] VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2_read_add;
wire [18:0] VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2;
VMStubs #("Tracklet") VMS_L4D3PHI2X2n4(
.data_in(VMR_L4D3_VMS_L4D3PHI2X2n4),
.enable(VMR_L4D3_VMS_L4D3PHI2X2n4_wr_en),
.number_out(VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2_number),
.read_add(VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2_read_add),
.data_out(VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X1n4;
wire VMR_L3D3_VMS_L3D3PHI2X1n4_wr_en;
wire [5:0] VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2_number;
wire [10:0] VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2_read_add;
wire [18:0] VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2;
VMStubs #("Tracklet") VMS_L3D3PHI2X1n4(
.data_in(VMR_L3D3_VMS_L3D3PHI2X1n4),
.enable(VMR_L3D3_VMS_L3D3PHI2X1n4_wr_en),
.number_out(VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2_number),
.read_add(VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2_read_add),
.data_out(VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X2n3;
wire VMR_L4D3_VMS_L4D3PHI3X2n3_wr_en;
wire [5:0] VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2_number;
wire [10:0] VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2_read_add;
wire [18:0] VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2;
VMStubs #("Tracklet") VMS_L4D3PHI3X2n3(
.data_in(VMR_L4D3_VMS_L4D3PHI3X2n3),
.enable(VMR_L4D3_VMS_L4D3PHI3X2n3_wr_en),
.number_out(VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2_number),
.read_add(VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2_read_add),
.data_out(VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X1n3;
wire VMR_L3D3_VMS_L3D3PHI3X1n3_wr_en;
wire [5:0] VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2_number;
wire [10:0] VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2_read_add;
wire [18:0] VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2;
VMStubs #("Tracklet") VMS_L3D3PHI3X1n3(
.data_in(VMR_L3D3_VMS_L3D3PHI3X1n3),
.enable(VMR_L3D3_VMS_L3D3PHI3X1n3_wr_en),
.number_out(VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2_number),
.read_add(VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2_read_add),
.data_out(VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X2n4;
wire VMR_L4D3_VMS_L4D3PHI3X2n4_wr_en;
wire [5:0] VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2_number;
wire [10:0] VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2_read_add;
wire [18:0] VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2;
VMStubs #("Tracklet") VMS_L4D3PHI3X2n4(
.data_in(VMR_L4D3_VMS_L4D3PHI3X2n4),
.enable(VMR_L4D3_VMS_L4D3PHI3X2n4_wr_en),
.number_out(VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2_number),
.read_add(VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2_read_add),
.data_out(VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X1n4;
wire VMR_L3D3_VMS_L3D3PHI3X1n4_wr_en;
wire [5:0] VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2_number;
wire [10:0] VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2_read_add;
wire [18:0] VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2;
VMStubs #("Tracklet") VMS_L3D3PHI3X1n4(
.data_in(VMR_L3D3_VMS_L3D3PHI3X1n4),
.enable(VMR_L3D3_VMS_L3D3PHI3X1n4_wr_en),
.number_out(VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2_number),
.read_add(VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2_read_add),
.data_out(VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI4X2n2;
wire VMR_L4D3_VMS_L4D3PHI4X2n2_wr_en;
wire [5:0] VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2_number;
wire [10:0] VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2_read_add;
wire [18:0] VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2;
VMStubs #("Tracklet") VMS_L4D3PHI4X2n2(
.data_in(VMR_L4D3_VMS_L4D3PHI4X2n2),
.enable(VMR_L4D3_VMS_L4D3PHI4X2n2_wr_en),
.number_out(VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2_number),
.read_add(VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2_read_add),
.data_out(VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X2n3;
wire VMR_L3D3_VMS_L3D3PHI1X2n3_wr_en;
wire [5:0] VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1_number;
wire [10:0] VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1_read_add;
wire [18:0] VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1;
VMStubs #("Tracklet") VMS_L3D3PHI1X2n3(
.data_in(VMR_L3D3_VMS_L3D3PHI1X2n3),
.enable(VMR_L3D3_VMS_L3D3PHI1X2n3_wr_en),
.number_out(VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1_number),
.read_add(VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1_read_add),
.data_out(VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI1X1n1;
wire VMR_L4D4_VMS_L4D4PHI1X1n1_wr_en;
wire [5:0] VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1_number;
wire [10:0] VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1_read_add;
wire [18:0] VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1;
VMStubs #("Tracklet") VMS_L4D4PHI1X1n1(
.data_in(VMR_L4D4_VMS_L4D4PHI1X1n1),
.enable(VMR_L4D4_VMS_L4D4PHI1X1n1_wr_en),
.number_out(VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1_number),
.read_add(VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1_read_add),
.data_out(VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X2n4;
wire VMR_L3D3_VMS_L3D3PHI1X2n4_wr_en;
wire [5:0] VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1_number;
wire [10:0] VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1_read_add;
wire [18:0] VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1;
VMStubs #("Tracklet") VMS_L3D3PHI1X2n4(
.data_in(VMR_L3D3_VMS_L3D3PHI1X2n4),
.enable(VMR_L3D3_VMS_L3D3PHI1X2n4_wr_en),
.number_out(VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1_number),
.read_add(VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1_read_add),
.data_out(VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X1n1;
wire VMR_L4D4_VMS_L4D4PHI2X1n1_wr_en;
wire [5:0] VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1_number;
wire [10:0] VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1_read_add;
wire [18:0] VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1;
VMStubs #("Tracklet") VMS_L4D4PHI2X1n1(
.data_in(VMR_L4D4_VMS_L4D4PHI2X1n1),
.enable(VMR_L4D4_VMS_L4D4PHI2X1n1_wr_en),
.number_out(VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1_number),
.read_add(VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1_read_add),
.data_out(VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X2n3;
wire VMR_L3D3_VMS_L3D3PHI2X2n3_wr_en;
wire [5:0] VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1_number;
wire [10:0] VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1_read_add;
wire [18:0] VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1;
VMStubs #("Tracklet") VMS_L3D3PHI2X2n3(
.data_in(VMR_L3D3_VMS_L3D3PHI2X2n3),
.enable(VMR_L3D3_VMS_L3D3PHI2X2n3_wr_en),
.number_out(VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1_number),
.read_add(VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1_read_add),
.data_out(VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X1n2;
wire VMR_L4D4_VMS_L4D4PHI2X1n2_wr_en;
wire [5:0] VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1_number;
wire [10:0] VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1_read_add;
wire [18:0] VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1;
VMStubs #("Tracklet") VMS_L4D4PHI2X1n2(
.data_in(VMR_L4D4_VMS_L4D4PHI2X1n2),
.enable(VMR_L4D4_VMS_L4D4PHI2X1n2_wr_en),
.number_out(VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1_number),
.read_add(VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1_read_add),
.data_out(VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X2n4;
wire VMR_L3D3_VMS_L3D3PHI2X2n4_wr_en;
wire [5:0] VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1_number;
wire [10:0] VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1_read_add;
wire [18:0] VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1;
VMStubs #("Tracklet") VMS_L3D3PHI2X2n4(
.data_in(VMR_L3D3_VMS_L3D3PHI2X2n4),
.enable(VMR_L3D3_VMS_L3D3PHI2X2n4_wr_en),
.number_out(VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1_number),
.read_add(VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1_read_add),
.data_out(VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X1n1;
wire VMR_L4D4_VMS_L4D4PHI3X1n1_wr_en;
wire [5:0] VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1_number;
wire [10:0] VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1_read_add;
wire [18:0] VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1;
VMStubs #("Tracklet") VMS_L4D4PHI3X1n1(
.data_in(VMR_L4D4_VMS_L4D4PHI3X1n1),
.enable(VMR_L4D4_VMS_L4D4PHI3X1n1_wr_en),
.number_out(VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1_number),
.read_add(VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1_read_add),
.data_out(VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X2n3;
wire VMR_L3D3_VMS_L3D3PHI3X2n3_wr_en;
wire [5:0] VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1_number;
wire [10:0] VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1_read_add;
wire [18:0] VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1;
VMStubs #("Tracklet") VMS_L3D3PHI3X2n3(
.data_in(VMR_L3D3_VMS_L3D3PHI3X2n3),
.enable(VMR_L3D3_VMS_L3D3PHI3X2n3_wr_en),
.number_out(VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1_number),
.read_add(VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1_read_add),
.data_out(VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X1n2;
wire VMR_L4D4_VMS_L4D4PHI3X1n2_wr_en;
wire [5:0] VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1_number;
wire [10:0] VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1_read_add;
wire [18:0] VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1;
VMStubs #("Tracklet") VMS_L4D4PHI3X1n2(
.data_in(VMR_L4D4_VMS_L4D4PHI3X1n2),
.enable(VMR_L4D4_VMS_L4D4PHI3X1n2_wr_en),
.number_out(VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1_number),
.read_add(VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1_read_add),
.data_out(VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X2n4;
wire VMR_L3D3_VMS_L3D3PHI3X2n4_wr_en;
wire [5:0] VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1_number;
wire [10:0] VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1_read_add;
wire [18:0] VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1;
VMStubs #("Tracklet") VMS_L3D3PHI3X2n4(
.data_in(VMR_L3D3_VMS_L3D3PHI3X2n4),
.enable(VMR_L3D3_VMS_L3D3PHI3X2n4_wr_en),
.number_out(VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1_number),
.read_add(VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1_read_add),
.data_out(VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI4X1n1;
wire VMR_L4D4_VMS_L4D4PHI4X1n1_wr_en;
wire [5:0] VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1_number;
wire [10:0] VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1_read_add;
wire [18:0] VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1;
VMStubs #("Tracklet") VMS_L4D4PHI4X1n1(
.data_in(VMR_L4D4_VMS_L4D4PHI4X1n1),
.enable(VMR_L4D4_VMS_L4D4PHI4X1n1_wr_en),
.number_out(VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1_number),
.read_add(VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1_read_add),
.data_out(VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X1n1;
wire VMR_L3D4_VMS_L3D4PHI1X1n1_wr_en;
wire [5:0] VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1_number;
wire [10:0] VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1_read_add;
wire [18:0] VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1;
VMStubs #("Tracklet") VMS_L3D4PHI1X1n1(
.data_in(VMR_L3D4_VMS_L3D4PHI1X1n1),
.enable(VMR_L3D4_VMS_L3D4PHI1X1n1_wr_en),
.number_out(VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1_number),
.read_add(VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1_read_add),
.data_out(VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI1X1n2;
wire VMR_L4D4_VMS_L4D4PHI1X1n2_wr_en;
wire [5:0] VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1_number;
wire [10:0] VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1_read_add;
wire [18:0] VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1;
VMStubs #("Tracklet") VMS_L4D4PHI1X1n2(
.data_in(VMR_L4D4_VMS_L4D4PHI1X1n2),
.enable(VMR_L4D4_VMS_L4D4PHI1X1n2_wr_en),
.number_out(VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1_number),
.read_add(VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1_read_add),
.data_out(VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X1n2;
wire VMR_L3D4_VMS_L3D4PHI1X1n2_wr_en;
wire [5:0] VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1_number;
wire [10:0] VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1_read_add;
wire [18:0] VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1;
VMStubs #("Tracklet") VMS_L3D4PHI1X1n2(
.data_in(VMR_L3D4_VMS_L3D4PHI1X1n2),
.enable(VMR_L3D4_VMS_L3D4PHI1X1n2_wr_en),
.number_out(VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1_number),
.read_add(VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1_read_add),
.data_out(VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X1n3;
wire VMR_L4D4_VMS_L4D4PHI2X1n3_wr_en;
wire [5:0] VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1_number;
wire [10:0] VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1_read_add;
wire [18:0] VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1;
VMStubs #("Tracklet") VMS_L4D4PHI2X1n3(
.data_in(VMR_L4D4_VMS_L4D4PHI2X1n3),
.enable(VMR_L4D4_VMS_L4D4PHI2X1n3_wr_en),
.number_out(VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1_number),
.read_add(VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1_read_add),
.data_out(VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X1n1;
wire VMR_L3D4_VMS_L3D4PHI2X1n1_wr_en;
wire [5:0] VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1_number;
wire [10:0] VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1_read_add;
wire [18:0] VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1;
VMStubs #("Tracklet") VMS_L3D4PHI2X1n1(
.data_in(VMR_L3D4_VMS_L3D4PHI2X1n1),
.enable(VMR_L3D4_VMS_L3D4PHI2X1n1_wr_en),
.number_out(VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1_number),
.read_add(VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1_read_add),
.data_out(VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X1n4;
wire VMR_L4D4_VMS_L4D4PHI2X1n4_wr_en;
wire [5:0] VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1_number;
wire [10:0] VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1_read_add;
wire [18:0] VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1;
VMStubs #("Tracklet") VMS_L4D4PHI2X1n4(
.data_in(VMR_L4D4_VMS_L4D4PHI2X1n4),
.enable(VMR_L4D4_VMS_L4D4PHI2X1n4_wr_en),
.number_out(VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1_number),
.read_add(VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1_read_add),
.data_out(VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X1n2;
wire VMR_L3D4_VMS_L3D4PHI2X1n2_wr_en;
wire [5:0] VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1_number;
wire [10:0] VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1_read_add;
wire [18:0] VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1;
VMStubs #("Tracklet") VMS_L3D4PHI2X1n2(
.data_in(VMR_L3D4_VMS_L3D4PHI2X1n2),
.enable(VMR_L3D4_VMS_L3D4PHI2X1n2_wr_en),
.number_out(VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1_number),
.read_add(VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1_read_add),
.data_out(VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X1n3;
wire VMR_L4D4_VMS_L4D4PHI3X1n3_wr_en;
wire [5:0] VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1_number;
wire [10:0] VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1_read_add;
wire [18:0] VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1;
VMStubs #("Tracklet") VMS_L4D4PHI3X1n3(
.data_in(VMR_L4D4_VMS_L4D4PHI3X1n3),
.enable(VMR_L4D4_VMS_L4D4PHI3X1n3_wr_en),
.number_out(VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1_number),
.read_add(VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1_read_add),
.data_out(VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X1n1;
wire VMR_L3D4_VMS_L3D4PHI3X1n1_wr_en;
wire [5:0] VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1_number;
wire [10:0] VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1_read_add;
wire [18:0] VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1;
VMStubs #("Tracklet") VMS_L3D4PHI3X1n1(
.data_in(VMR_L3D4_VMS_L3D4PHI3X1n1),
.enable(VMR_L3D4_VMS_L3D4PHI3X1n1_wr_en),
.number_out(VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1_number),
.read_add(VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1_read_add),
.data_out(VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X1n4;
wire VMR_L4D4_VMS_L4D4PHI3X1n4_wr_en;
wire [5:0] VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1_number;
wire [10:0] VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1_read_add;
wire [18:0] VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1;
VMStubs #("Tracklet") VMS_L4D4PHI3X1n4(
.data_in(VMR_L4D4_VMS_L4D4PHI3X1n4),
.enable(VMR_L4D4_VMS_L4D4PHI3X1n4_wr_en),
.number_out(VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1_number),
.read_add(VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1_read_add),
.data_out(VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X1n2;
wire VMR_L3D4_VMS_L3D4PHI3X1n2_wr_en;
wire [5:0] VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_number;
wire [10:0] VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_read_add;
wire [18:0] VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1;
VMStubs #("Tracklet") VMS_L3D4PHI3X1n2(
.data_in(VMR_L3D4_VMS_L3D4PHI3X1n2),
.enable(VMR_L3D4_VMS_L3D4PHI3X1n2_wr_en),
.number_out(VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_number),
.read_add(VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_read_add),
.data_out(VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI4X1n2;
wire VMR_L4D4_VMS_L4D4PHI4X1n2_wr_en;
wire [5:0] VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_number;
wire [10:0] VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_read_add;
wire [18:0] VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1;
VMStubs #("Tracklet") VMS_L4D4PHI4X1n2(
.data_in(VMR_L4D4_VMS_L4D4PHI4X1n2),
.enable(VMR_L4D4_VMS_L4D4PHI4X1n2_wr_en),
.number_out(VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_number),
.read_add(VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_read_add),
.data_out(VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X1n3;
wire VMR_L3D4_VMS_L3D4PHI1X1n3_wr_en;
wire [5:0] VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2_number;
wire [10:0] VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2_read_add;
wire [18:0] VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2;
VMStubs #("Tracklet") VMS_L3D4PHI1X1n3(
.data_in(VMR_L3D4_VMS_L3D4PHI1X1n3),
.enable(VMR_L3D4_VMS_L3D4PHI1X1n3_wr_en),
.number_out(VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2_number),
.read_add(VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2_read_add),
.data_out(VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI1X2n1;
wire VMR_L4D4_VMS_L4D4PHI1X2n1_wr_en;
wire [5:0] VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2_number;
wire [10:0] VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2_read_add;
wire [18:0] VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2;
VMStubs #("Tracklet") VMS_L4D4PHI1X2n1(
.data_in(VMR_L4D4_VMS_L4D4PHI1X2n1),
.enable(VMR_L4D4_VMS_L4D4PHI1X2n1_wr_en),
.number_out(VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2_number),
.read_add(VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2_read_add),
.data_out(VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X1n4;
wire VMR_L3D4_VMS_L3D4PHI1X1n4_wr_en;
wire [5:0] VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2_number;
wire [10:0] VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2_read_add;
wire [18:0] VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2;
VMStubs #("Tracklet") VMS_L3D4PHI1X1n4(
.data_in(VMR_L3D4_VMS_L3D4PHI1X1n4),
.enable(VMR_L3D4_VMS_L3D4PHI1X1n4_wr_en),
.number_out(VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2_number),
.read_add(VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2_read_add),
.data_out(VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X2n1;
wire VMR_L4D4_VMS_L4D4PHI2X2n1_wr_en;
wire [5:0] VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2_number;
wire [10:0] VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2_read_add;
wire [18:0] VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2;
VMStubs #("Tracklet") VMS_L4D4PHI2X2n1(
.data_in(VMR_L4D4_VMS_L4D4PHI2X2n1),
.enable(VMR_L4D4_VMS_L4D4PHI2X2n1_wr_en),
.number_out(VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2_number),
.read_add(VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2_read_add),
.data_out(VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X1n3;
wire VMR_L3D4_VMS_L3D4PHI2X1n3_wr_en;
wire [5:0] VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2_number;
wire [10:0] VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2_read_add;
wire [18:0] VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2;
VMStubs #("Tracklet") VMS_L3D4PHI2X1n3(
.data_in(VMR_L3D4_VMS_L3D4PHI2X1n3),
.enable(VMR_L3D4_VMS_L3D4PHI2X1n3_wr_en),
.number_out(VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2_number),
.read_add(VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2_read_add),
.data_out(VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X2n2;
wire VMR_L4D4_VMS_L4D4PHI2X2n2_wr_en;
wire [5:0] VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2_number;
wire [10:0] VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2_read_add;
wire [18:0] VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2;
VMStubs #("Tracklet") VMS_L4D4PHI2X2n2(
.data_in(VMR_L4D4_VMS_L4D4PHI2X2n2),
.enable(VMR_L4D4_VMS_L4D4PHI2X2n2_wr_en),
.number_out(VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2_number),
.read_add(VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2_read_add),
.data_out(VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X1n4;
wire VMR_L3D4_VMS_L3D4PHI2X1n4_wr_en;
wire [5:0] VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2_number;
wire [10:0] VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2_read_add;
wire [18:0] VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2;
VMStubs #("Tracklet") VMS_L3D4PHI2X1n4(
.data_in(VMR_L3D4_VMS_L3D4PHI2X1n4),
.enable(VMR_L3D4_VMS_L3D4PHI2X1n4_wr_en),
.number_out(VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2_number),
.read_add(VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2_read_add),
.data_out(VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X2n1;
wire VMR_L4D4_VMS_L4D4PHI3X2n1_wr_en;
wire [5:0] VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2_number;
wire [10:0] VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2_read_add;
wire [18:0] VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2;
VMStubs #("Tracklet") VMS_L4D4PHI3X2n1(
.data_in(VMR_L4D4_VMS_L4D4PHI3X2n1),
.enable(VMR_L4D4_VMS_L4D4PHI3X2n1_wr_en),
.number_out(VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2_number),
.read_add(VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2_read_add),
.data_out(VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X1n3;
wire VMR_L3D4_VMS_L3D4PHI3X1n3_wr_en;
wire [5:0] VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2_number;
wire [10:0] VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2_read_add;
wire [18:0] VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2;
VMStubs #("Tracklet") VMS_L3D4PHI3X1n3(
.data_in(VMR_L3D4_VMS_L3D4PHI3X1n3),
.enable(VMR_L3D4_VMS_L3D4PHI3X1n3_wr_en),
.number_out(VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2_number),
.read_add(VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2_read_add),
.data_out(VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X2n2;
wire VMR_L4D4_VMS_L4D4PHI3X2n2_wr_en;
wire [5:0] VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2_number;
wire [10:0] VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2_read_add;
wire [18:0] VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2;
VMStubs #("Tracklet") VMS_L4D4PHI3X2n2(
.data_in(VMR_L4D4_VMS_L4D4PHI3X2n2),
.enable(VMR_L4D4_VMS_L4D4PHI3X2n2_wr_en),
.number_out(VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2_number),
.read_add(VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2_read_add),
.data_out(VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X1n4;
wire VMR_L3D4_VMS_L3D4PHI3X1n4_wr_en;
wire [5:0] VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2_number;
wire [10:0] VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2_read_add;
wire [18:0] VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2;
VMStubs #("Tracklet") VMS_L3D4PHI3X1n4(
.data_in(VMR_L3D4_VMS_L3D4PHI3X1n4),
.enable(VMR_L3D4_VMS_L3D4PHI3X1n4_wr_en),
.number_out(VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2_number),
.read_add(VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2_read_add),
.data_out(VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI4X2n1;
wire VMR_L4D4_VMS_L4D4PHI4X2n1_wr_en;
wire [5:0] VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2_number;
wire [10:0] VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2_read_add;
wire [18:0] VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2;
VMStubs #("Tracklet") VMS_L4D4PHI4X2n1(
.data_in(VMR_L4D4_VMS_L4D4PHI4X2n1),
.enable(VMR_L4D4_VMS_L4D4PHI4X2n1_wr_en),
.number_out(VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2_number),
.read_add(VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2_read_add),
.data_out(VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X2n1;
wire VMR_L3D4_VMS_L3D4PHI1X2n1_wr_en;
wire [5:0] VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2_number;
wire [10:0] VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2_read_add;
wire [18:0] VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2;
VMStubs #("Tracklet") VMS_L3D4PHI1X2n1(
.data_in(VMR_L3D4_VMS_L3D4PHI1X2n1),
.enable(VMR_L3D4_VMS_L3D4PHI1X2n1_wr_en),
.number_out(VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2_number),
.read_add(VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2_read_add),
.data_out(VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI1X2n2;
wire VMR_L4D4_VMS_L4D4PHI1X2n2_wr_en;
wire [5:0] VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2_number;
wire [10:0] VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2_read_add;
wire [18:0] VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2;
VMStubs #("Tracklet") VMS_L4D4PHI1X2n2(
.data_in(VMR_L4D4_VMS_L4D4PHI1X2n2),
.enable(VMR_L4D4_VMS_L4D4PHI1X2n2_wr_en),
.number_out(VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2_number),
.read_add(VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2_read_add),
.data_out(VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X2n2;
wire VMR_L3D4_VMS_L3D4PHI1X2n2_wr_en;
wire [5:0] VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2_number;
wire [10:0] VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2_read_add;
wire [18:0] VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2;
VMStubs #("Tracklet") VMS_L3D4PHI1X2n2(
.data_in(VMR_L3D4_VMS_L3D4PHI1X2n2),
.enable(VMR_L3D4_VMS_L3D4PHI1X2n2_wr_en),
.number_out(VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2_number),
.read_add(VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2_read_add),
.data_out(VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X2n3;
wire VMR_L4D4_VMS_L4D4PHI2X2n3_wr_en;
wire [5:0] VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2_number;
wire [10:0] VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2_read_add;
wire [18:0] VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2;
VMStubs #("Tracklet") VMS_L4D4PHI2X2n3(
.data_in(VMR_L4D4_VMS_L4D4PHI2X2n3),
.enable(VMR_L4D4_VMS_L4D4PHI2X2n3_wr_en),
.number_out(VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2_number),
.read_add(VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2_read_add),
.data_out(VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X2n1;
wire VMR_L3D4_VMS_L3D4PHI2X2n1_wr_en;
wire [5:0] VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2_number;
wire [10:0] VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2_read_add;
wire [18:0] VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2;
VMStubs #("Tracklet") VMS_L3D4PHI2X2n1(
.data_in(VMR_L3D4_VMS_L3D4PHI2X2n1),
.enable(VMR_L3D4_VMS_L3D4PHI2X2n1_wr_en),
.number_out(VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2_number),
.read_add(VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2_read_add),
.data_out(VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X2n4;
wire VMR_L4D4_VMS_L4D4PHI2X2n4_wr_en;
wire [5:0] VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2_number;
wire [10:0] VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2_read_add;
wire [18:0] VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2;
VMStubs #("Tracklet") VMS_L4D4PHI2X2n4(
.data_in(VMR_L4D4_VMS_L4D4PHI2X2n4),
.enable(VMR_L4D4_VMS_L4D4PHI2X2n4_wr_en),
.number_out(VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2_number),
.read_add(VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2_read_add),
.data_out(VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X2n2;
wire VMR_L3D4_VMS_L3D4PHI2X2n2_wr_en;
wire [5:0] VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2_number;
wire [10:0] VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2_read_add;
wire [18:0] VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2;
VMStubs #("Tracklet") VMS_L3D4PHI2X2n2(
.data_in(VMR_L3D4_VMS_L3D4PHI2X2n2),
.enable(VMR_L3D4_VMS_L3D4PHI2X2n2_wr_en),
.number_out(VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2_number),
.read_add(VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2_read_add),
.data_out(VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X2n3;
wire VMR_L4D4_VMS_L4D4PHI3X2n3_wr_en;
wire [5:0] VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2_number;
wire [10:0] VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2_read_add;
wire [18:0] VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2;
VMStubs #("Tracklet") VMS_L4D4PHI3X2n3(
.data_in(VMR_L4D4_VMS_L4D4PHI3X2n3),
.enable(VMR_L4D4_VMS_L4D4PHI3X2n3_wr_en),
.number_out(VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2_number),
.read_add(VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2_read_add),
.data_out(VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X2n1;
wire VMR_L3D4_VMS_L3D4PHI3X2n1_wr_en;
wire [5:0] VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2_number;
wire [10:0] VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2_read_add;
wire [18:0] VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2;
VMStubs #("Tracklet") VMS_L3D4PHI3X2n1(
.data_in(VMR_L3D4_VMS_L3D4PHI3X2n1),
.enable(VMR_L3D4_VMS_L3D4PHI3X2n1_wr_en),
.number_out(VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2_number),
.read_add(VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2_read_add),
.data_out(VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X2n4;
wire VMR_L4D4_VMS_L4D4PHI3X2n4_wr_en;
wire [5:0] VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2_number;
wire [10:0] VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2_read_add;
wire [18:0] VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2;
VMStubs #("Tracklet") VMS_L4D4PHI3X2n4(
.data_in(VMR_L4D4_VMS_L4D4PHI3X2n4),
.enable(VMR_L4D4_VMS_L4D4PHI3X2n4_wr_en),
.number_out(VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2_number),
.read_add(VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2_read_add),
.data_out(VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X2n2;
wire VMR_L3D4_VMS_L3D4PHI3X2n2_wr_en;
wire [5:0] VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_number;
wire [10:0] VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_read_add;
wire [18:0] VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2;
VMStubs #("Tracklet") VMS_L3D4PHI3X2n2(
.data_in(VMR_L3D4_VMS_L3D4PHI3X2n2),
.enable(VMR_L3D4_VMS_L3D4PHI3X2n2_wr_en),
.number_out(VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_number),
.read_add(VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_read_add),
.data_out(VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI4X2n2;
wire VMR_L4D4_VMS_L4D4PHI4X2n2_wr_en;
wire [5:0] VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_number;
wire [10:0] VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_read_add;
wire [18:0] VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2;
VMStubs #("Tracklet") VMS_L4D4PHI4X2n2(
.data_in(VMR_L4D4_VMS_L4D4PHI4X2n2),
.enable(VMR_L4D4_VMS_L4D4PHI4X2n2_wr_en),
.number_out(VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_number),
.read_add(VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_read_add),
.data_out(VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X1n1;
wire VMR_L5D3_VMS_L5D3PHI1X1n1_wr_en;
wire [5:0] VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_number;
wire [10:0] VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_read_add;
wire [18:0] VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1;
VMStubs #("Tracklet") VMS_L5D3PHI1X1n1(
.data_in(VMR_L5D3_VMS_L5D3PHI1X1n1),
.enable(VMR_L5D3_VMS_L5D3PHI1X1n1_wr_en),
.number_out(VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_number),
.read_add(VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_read_add),
.data_out(VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI1X1n1;
wire VMR_L6D3_VMS_L6D3PHI1X1n1_wr_en;
wire [5:0] VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_number;
wire [10:0] VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_read_add;
wire [18:0] VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1;
VMStubs #("Tracklet") VMS_L6D3PHI1X1n1(
.data_in(VMR_L6D3_VMS_L6D3PHI1X1n1),
.enable(VMR_L6D3_VMS_L6D3PHI1X1n1_wr_en),
.number_out(VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_number),
.read_add(VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_read_add),
.data_out(VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X1n2;
wire VMR_L5D3_VMS_L5D3PHI1X1n2_wr_en;
wire [5:0] VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1_number;
wire [10:0] VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1_read_add;
wire [18:0] VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1;
VMStubs #("Tracklet") VMS_L5D3PHI1X1n2(
.data_in(VMR_L5D3_VMS_L5D3PHI1X1n2),
.enable(VMR_L5D3_VMS_L5D3PHI1X1n2_wr_en),
.number_out(VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1_number),
.read_add(VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1_read_add),
.data_out(VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X1n1;
wire VMR_L6D3_VMS_L6D3PHI2X1n1_wr_en;
wire [5:0] VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1_number;
wire [10:0] VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1_read_add;
wire [18:0] VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1;
VMStubs #("Tracklet") VMS_L6D3PHI2X1n1(
.data_in(VMR_L6D3_VMS_L6D3PHI2X1n1),
.enable(VMR_L6D3_VMS_L6D3PHI2X1n1_wr_en),
.number_out(VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1_number),
.read_add(VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1_read_add),
.data_out(VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X1n1;
wire VMR_L5D3_VMS_L5D3PHI2X1n1_wr_en;
wire [5:0] VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1_number;
wire [10:0] VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1_read_add;
wire [18:0] VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1;
VMStubs #("Tracklet") VMS_L5D3PHI2X1n1(
.data_in(VMR_L5D3_VMS_L5D3PHI2X1n1),
.enable(VMR_L5D3_VMS_L5D3PHI2X1n1_wr_en),
.number_out(VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1_number),
.read_add(VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1_read_add),
.data_out(VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X1n2;
wire VMR_L6D3_VMS_L6D3PHI2X1n2_wr_en;
wire [5:0] VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1_number;
wire [10:0] VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1_read_add;
wire [18:0] VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1;
VMStubs #("Tracklet") VMS_L6D3PHI2X1n2(
.data_in(VMR_L6D3_VMS_L6D3PHI2X1n2),
.enable(VMR_L6D3_VMS_L6D3PHI2X1n2_wr_en),
.number_out(VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1_number),
.read_add(VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1_read_add),
.data_out(VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X1n2;
wire VMR_L5D3_VMS_L5D3PHI2X1n2_wr_en;
wire [5:0] VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1_number;
wire [10:0] VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1_read_add;
wire [18:0] VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1;
VMStubs #("Tracklet") VMS_L5D3PHI2X1n2(
.data_in(VMR_L5D3_VMS_L5D3PHI2X1n2),
.enable(VMR_L5D3_VMS_L5D3PHI2X1n2_wr_en),
.number_out(VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1_number),
.read_add(VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1_read_add),
.data_out(VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X1n1;
wire VMR_L6D3_VMS_L6D3PHI3X1n1_wr_en;
wire [5:0] VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1_number;
wire [10:0] VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1_read_add;
wire [18:0] VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1;
VMStubs #("Tracklet") VMS_L6D3PHI3X1n1(
.data_in(VMR_L6D3_VMS_L6D3PHI3X1n1),
.enable(VMR_L6D3_VMS_L6D3PHI3X1n1_wr_en),
.number_out(VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1_number),
.read_add(VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1_read_add),
.data_out(VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X1n1;
wire VMR_L5D3_VMS_L5D3PHI3X1n1_wr_en;
wire [5:0] VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1_number;
wire [10:0] VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1_read_add;
wire [18:0] VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1;
VMStubs #("Tracklet") VMS_L5D3PHI3X1n1(
.data_in(VMR_L5D3_VMS_L5D3PHI3X1n1),
.enable(VMR_L5D3_VMS_L5D3PHI3X1n1_wr_en),
.number_out(VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1_number),
.read_add(VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1_read_add),
.data_out(VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X1n2;
wire VMR_L6D3_VMS_L6D3PHI3X1n2_wr_en;
wire [5:0] VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1_number;
wire [10:0] VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1_read_add;
wire [18:0] VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1;
VMStubs #("Tracklet") VMS_L6D3PHI3X1n2(
.data_in(VMR_L6D3_VMS_L6D3PHI3X1n2),
.enable(VMR_L6D3_VMS_L6D3PHI3X1n2_wr_en),
.number_out(VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1_number),
.read_add(VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1_read_add),
.data_out(VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X1n2;
wire VMR_L5D3_VMS_L5D3PHI3X1n2_wr_en;
wire [5:0] VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1_number;
wire [10:0] VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1_read_add;
wire [18:0] VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1;
VMStubs #("Tracklet") VMS_L5D3PHI3X1n2(
.data_in(VMR_L5D3_VMS_L5D3PHI3X1n2),
.enable(VMR_L5D3_VMS_L5D3PHI3X1n2_wr_en),
.number_out(VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1_number),
.read_add(VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1_read_add),
.data_out(VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI4X1n1;
wire VMR_L6D3_VMS_L6D3PHI4X1n1_wr_en;
wire [5:0] VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1_number;
wire [10:0] VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1_read_add;
wire [18:0] VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1;
VMStubs #("Tracklet") VMS_L6D3PHI4X1n1(
.data_in(VMR_L6D3_VMS_L6D3PHI4X1n1),
.enable(VMR_L6D3_VMS_L6D3PHI4X1n1_wr_en),
.number_out(VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1_number),
.read_add(VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1_read_add),
.data_out(VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X1n3;
wire VMR_L5D3_VMS_L5D3PHI1X1n3_wr_en;
wire [5:0] VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2_number;
wire [10:0] VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2_read_add;
wire [18:0] VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2;
VMStubs #("Tracklet") VMS_L5D3PHI1X1n3(
.data_in(VMR_L5D3_VMS_L5D3PHI1X1n3),
.enable(VMR_L5D3_VMS_L5D3PHI1X1n3_wr_en),
.number_out(VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2_number),
.read_add(VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2_read_add),
.data_out(VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI1X2n1;
wire VMR_L6D3_VMS_L6D3PHI1X2n1_wr_en;
wire [5:0] VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2_number;
wire [10:0] VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2_read_add;
wire [18:0] VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2;
VMStubs #("Tracklet") VMS_L6D3PHI1X2n1(
.data_in(VMR_L6D3_VMS_L6D3PHI1X2n1),
.enable(VMR_L6D3_VMS_L6D3PHI1X2n1_wr_en),
.number_out(VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2_number),
.read_add(VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2_read_add),
.data_out(VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X1n4;
wire VMR_L5D3_VMS_L5D3PHI1X1n4_wr_en;
wire [5:0] VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2_number;
wire [10:0] VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2_read_add;
wire [18:0] VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2;
VMStubs #("Tracklet") VMS_L5D3PHI1X1n4(
.data_in(VMR_L5D3_VMS_L5D3PHI1X1n4),
.enable(VMR_L5D3_VMS_L5D3PHI1X1n4_wr_en),
.number_out(VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2_number),
.read_add(VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2_read_add),
.data_out(VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X2n1;
wire VMR_L6D3_VMS_L6D3PHI2X2n1_wr_en;
wire [5:0] VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2_number;
wire [10:0] VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2_read_add;
wire [18:0] VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2;
VMStubs #("Tracklet") VMS_L6D3PHI2X2n1(
.data_in(VMR_L6D3_VMS_L6D3PHI2X2n1),
.enable(VMR_L6D3_VMS_L6D3PHI2X2n1_wr_en),
.number_out(VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2_number),
.read_add(VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2_read_add),
.data_out(VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X1n3;
wire VMR_L5D3_VMS_L5D3PHI2X1n3_wr_en;
wire [5:0] VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2_number;
wire [10:0] VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2_read_add;
wire [18:0] VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2;
VMStubs #("Tracklet") VMS_L5D3PHI2X1n3(
.data_in(VMR_L5D3_VMS_L5D3PHI2X1n3),
.enable(VMR_L5D3_VMS_L5D3PHI2X1n3_wr_en),
.number_out(VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2_number),
.read_add(VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2_read_add),
.data_out(VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X2n2;
wire VMR_L6D3_VMS_L6D3PHI2X2n2_wr_en;
wire [5:0] VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2_number;
wire [10:0] VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2_read_add;
wire [18:0] VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2;
VMStubs #("Tracklet") VMS_L6D3PHI2X2n2(
.data_in(VMR_L6D3_VMS_L6D3PHI2X2n2),
.enable(VMR_L6D3_VMS_L6D3PHI2X2n2_wr_en),
.number_out(VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2_number),
.read_add(VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2_read_add),
.data_out(VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X1n4;
wire VMR_L5D3_VMS_L5D3PHI2X1n4_wr_en;
wire [5:0] VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2_number;
wire [10:0] VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2_read_add;
wire [18:0] VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2;
VMStubs #("Tracklet") VMS_L5D3PHI2X1n4(
.data_in(VMR_L5D3_VMS_L5D3PHI2X1n4),
.enable(VMR_L5D3_VMS_L5D3PHI2X1n4_wr_en),
.number_out(VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2_number),
.read_add(VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2_read_add),
.data_out(VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X2n1;
wire VMR_L6D3_VMS_L6D3PHI3X2n1_wr_en;
wire [5:0] VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2_number;
wire [10:0] VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2_read_add;
wire [18:0] VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2;
VMStubs #("Tracklet") VMS_L6D3PHI3X2n1(
.data_in(VMR_L6D3_VMS_L6D3PHI3X2n1),
.enable(VMR_L6D3_VMS_L6D3PHI3X2n1_wr_en),
.number_out(VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2_number),
.read_add(VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2_read_add),
.data_out(VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X1n3;
wire VMR_L5D3_VMS_L5D3PHI3X1n3_wr_en;
wire [5:0] VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2_number;
wire [10:0] VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2_read_add;
wire [18:0] VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2;
VMStubs #("Tracklet") VMS_L5D3PHI3X1n3(
.data_in(VMR_L5D3_VMS_L5D3PHI3X1n3),
.enable(VMR_L5D3_VMS_L5D3PHI3X1n3_wr_en),
.number_out(VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2_number),
.read_add(VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2_read_add),
.data_out(VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X2n2;
wire VMR_L6D3_VMS_L6D3PHI3X2n2_wr_en;
wire [5:0] VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2_number;
wire [10:0] VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2_read_add;
wire [18:0] VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2;
VMStubs #("Tracklet") VMS_L6D3PHI3X2n2(
.data_in(VMR_L6D3_VMS_L6D3PHI3X2n2),
.enable(VMR_L6D3_VMS_L6D3PHI3X2n2_wr_en),
.number_out(VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2_number),
.read_add(VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2_read_add),
.data_out(VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X1n4;
wire VMR_L5D3_VMS_L5D3PHI3X1n4_wr_en;
wire [5:0] VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2_number;
wire [10:0] VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2_read_add;
wire [18:0] VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2;
VMStubs #("Tracklet") VMS_L5D3PHI3X1n4(
.data_in(VMR_L5D3_VMS_L5D3PHI3X1n4),
.enable(VMR_L5D3_VMS_L5D3PHI3X1n4_wr_en),
.number_out(VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2_number),
.read_add(VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2_read_add),
.data_out(VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI4X2n1;
wire VMR_L6D3_VMS_L6D3PHI4X2n1_wr_en;
wire [5:0] VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2_number;
wire [10:0] VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2_read_add;
wire [18:0] VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2;
VMStubs #("Tracklet") VMS_L6D3PHI4X2n1(
.data_in(VMR_L6D3_VMS_L6D3PHI4X2n1),
.enable(VMR_L6D3_VMS_L6D3PHI4X2n1_wr_en),
.number_out(VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2_number),
.read_add(VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2_read_add),
.data_out(VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X2n1;
wire VMR_L5D3_VMS_L5D3PHI1X2n1_wr_en;
wire [5:0] VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2_number;
wire [10:0] VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2_read_add;
wire [18:0] VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2;
VMStubs #("Tracklet") VMS_L5D3PHI1X2n1(
.data_in(VMR_L5D3_VMS_L5D3PHI1X2n1),
.enable(VMR_L5D3_VMS_L5D3PHI1X2n1_wr_en),
.number_out(VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2_number),
.read_add(VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2_read_add),
.data_out(VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI1X2n2;
wire VMR_L6D3_VMS_L6D3PHI1X2n2_wr_en;
wire [5:0] VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2_number;
wire [10:0] VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2_read_add;
wire [18:0] VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2;
VMStubs #("Tracklet") VMS_L6D3PHI1X2n2(
.data_in(VMR_L6D3_VMS_L6D3PHI1X2n2),
.enable(VMR_L6D3_VMS_L6D3PHI1X2n2_wr_en),
.number_out(VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2_number),
.read_add(VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2_read_add),
.data_out(VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X2n2;
wire VMR_L5D3_VMS_L5D3PHI1X2n2_wr_en;
wire [5:0] VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2_number;
wire [10:0] VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2_read_add;
wire [18:0] VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2;
VMStubs #("Tracklet") VMS_L5D3PHI1X2n2(
.data_in(VMR_L5D3_VMS_L5D3PHI1X2n2),
.enable(VMR_L5D3_VMS_L5D3PHI1X2n2_wr_en),
.number_out(VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2_number),
.read_add(VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2_read_add),
.data_out(VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X2n3;
wire VMR_L6D3_VMS_L6D3PHI2X2n3_wr_en;
wire [5:0] VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2_number;
wire [10:0] VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2_read_add;
wire [18:0] VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2;
VMStubs #("Tracklet") VMS_L6D3PHI2X2n3(
.data_in(VMR_L6D3_VMS_L6D3PHI2X2n3),
.enable(VMR_L6D3_VMS_L6D3PHI2X2n3_wr_en),
.number_out(VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2_number),
.read_add(VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2_read_add),
.data_out(VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X2n1;
wire VMR_L5D3_VMS_L5D3PHI2X2n1_wr_en;
wire [5:0] VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2_number;
wire [10:0] VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2_read_add;
wire [18:0] VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2;
VMStubs #("Tracklet") VMS_L5D3PHI2X2n1(
.data_in(VMR_L5D3_VMS_L5D3PHI2X2n1),
.enable(VMR_L5D3_VMS_L5D3PHI2X2n1_wr_en),
.number_out(VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2_number),
.read_add(VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2_read_add),
.data_out(VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X2n4;
wire VMR_L6D3_VMS_L6D3PHI2X2n4_wr_en;
wire [5:0] VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2_number;
wire [10:0] VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2_read_add;
wire [18:0] VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2;
VMStubs #("Tracklet") VMS_L6D3PHI2X2n4(
.data_in(VMR_L6D3_VMS_L6D3PHI2X2n4),
.enable(VMR_L6D3_VMS_L6D3PHI2X2n4_wr_en),
.number_out(VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2_number),
.read_add(VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2_read_add),
.data_out(VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X2n2;
wire VMR_L5D3_VMS_L5D3PHI2X2n2_wr_en;
wire [5:0] VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2_number;
wire [10:0] VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2_read_add;
wire [18:0] VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2;
VMStubs #("Tracklet") VMS_L5D3PHI2X2n2(
.data_in(VMR_L5D3_VMS_L5D3PHI2X2n2),
.enable(VMR_L5D3_VMS_L5D3PHI2X2n2_wr_en),
.number_out(VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2_number),
.read_add(VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2_read_add),
.data_out(VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X2n3;
wire VMR_L6D3_VMS_L6D3PHI3X2n3_wr_en;
wire [5:0] VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2_number;
wire [10:0] VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2_read_add;
wire [18:0] VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2;
VMStubs #("Tracklet") VMS_L6D3PHI3X2n3(
.data_in(VMR_L6D3_VMS_L6D3PHI3X2n3),
.enable(VMR_L6D3_VMS_L6D3PHI3X2n3_wr_en),
.number_out(VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2_number),
.read_add(VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2_read_add),
.data_out(VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X2n1;
wire VMR_L5D3_VMS_L5D3PHI3X2n1_wr_en;
wire [5:0] VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2_number;
wire [10:0] VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2_read_add;
wire [18:0] VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2;
VMStubs #("Tracklet") VMS_L5D3PHI3X2n1(
.data_in(VMR_L5D3_VMS_L5D3PHI3X2n1),
.enable(VMR_L5D3_VMS_L5D3PHI3X2n1_wr_en),
.number_out(VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2_number),
.read_add(VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2_read_add),
.data_out(VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X2n4;
wire VMR_L6D3_VMS_L6D3PHI3X2n4_wr_en;
wire [5:0] VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2_number;
wire [10:0] VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2_read_add;
wire [18:0] VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2;
VMStubs #("Tracklet") VMS_L6D3PHI3X2n4(
.data_in(VMR_L6D3_VMS_L6D3PHI3X2n4),
.enable(VMR_L6D3_VMS_L6D3PHI3X2n4_wr_en),
.number_out(VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2_number),
.read_add(VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2_read_add),
.data_out(VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X2n2;
wire VMR_L5D3_VMS_L5D3PHI3X2n2_wr_en;
wire [5:0] VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_number;
wire [10:0] VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_read_add;
wire [18:0] VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2;
VMStubs #("Tracklet") VMS_L5D3PHI3X2n2(
.data_in(VMR_L5D3_VMS_L5D3PHI3X2n2),
.enable(VMR_L5D3_VMS_L5D3PHI3X2n2_wr_en),
.number_out(VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_number),
.read_add(VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_read_add),
.data_out(VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI4X2n2;
wire VMR_L6D3_VMS_L6D3PHI4X2n2_wr_en;
wire [5:0] VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_number;
wire [10:0] VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_read_add;
wire [18:0] VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2;
VMStubs #("Tracklet") VMS_L6D3PHI4X2n2(
.data_in(VMR_L6D3_VMS_L6D3PHI4X2n2),
.enable(VMR_L6D3_VMS_L6D3PHI4X2n2_wr_en),
.number_out(VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_number),
.read_add(VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_read_add),
.data_out(VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X2n3;
wire VMR_L5D3_VMS_L5D3PHI1X2n3_wr_en;
wire [5:0] VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1_number;
wire [10:0] VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1_read_add;
wire [18:0] VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1;
VMStubs #("Tracklet") VMS_L5D3PHI1X2n3(
.data_in(VMR_L5D3_VMS_L5D3PHI1X2n3),
.enable(VMR_L5D3_VMS_L5D3PHI1X2n3_wr_en),
.number_out(VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1_number),
.read_add(VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1_read_add),
.data_out(VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI1X1n1;
wire VMR_L6D4_VMS_L6D4PHI1X1n1_wr_en;
wire [5:0] VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1_number;
wire [10:0] VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1_read_add;
wire [18:0] VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1;
VMStubs #("Tracklet") VMS_L6D4PHI1X1n1(
.data_in(VMR_L6D4_VMS_L6D4PHI1X1n1),
.enable(VMR_L6D4_VMS_L6D4PHI1X1n1_wr_en),
.number_out(VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1_number),
.read_add(VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1_read_add),
.data_out(VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X2n4;
wire VMR_L5D3_VMS_L5D3PHI1X2n4_wr_en;
wire [5:0] VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1_number;
wire [10:0] VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1_read_add;
wire [18:0] VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1;
VMStubs #("Tracklet") VMS_L5D3PHI1X2n4(
.data_in(VMR_L5D3_VMS_L5D3PHI1X2n4),
.enable(VMR_L5D3_VMS_L5D3PHI1X2n4_wr_en),
.number_out(VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1_number),
.read_add(VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1_read_add),
.data_out(VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X1n1;
wire VMR_L6D4_VMS_L6D4PHI2X1n1_wr_en;
wire [5:0] VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1_number;
wire [10:0] VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1_read_add;
wire [18:0] VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1;
VMStubs #("Tracklet") VMS_L6D4PHI2X1n1(
.data_in(VMR_L6D4_VMS_L6D4PHI2X1n1),
.enable(VMR_L6D4_VMS_L6D4PHI2X1n1_wr_en),
.number_out(VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1_number),
.read_add(VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1_read_add),
.data_out(VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X2n3;
wire VMR_L5D3_VMS_L5D3PHI2X2n3_wr_en;
wire [5:0] VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1_number;
wire [10:0] VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1_read_add;
wire [18:0] VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1;
VMStubs #("Tracklet") VMS_L5D3PHI2X2n3(
.data_in(VMR_L5D3_VMS_L5D3PHI2X2n3),
.enable(VMR_L5D3_VMS_L5D3PHI2X2n3_wr_en),
.number_out(VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1_number),
.read_add(VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1_read_add),
.data_out(VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X1n2;
wire VMR_L6D4_VMS_L6D4PHI2X1n2_wr_en;
wire [5:0] VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1_number;
wire [10:0] VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1_read_add;
wire [18:0] VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1;
VMStubs #("Tracklet") VMS_L6D4PHI2X1n2(
.data_in(VMR_L6D4_VMS_L6D4PHI2X1n2),
.enable(VMR_L6D4_VMS_L6D4PHI2X1n2_wr_en),
.number_out(VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1_number),
.read_add(VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1_read_add),
.data_out(VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X2n4;
wire VMR_L5D3_VMS_L5D3PHI2X2n4_wr_en;
wire [5:0] VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1_number;
wire [10:0] VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1_read_add;
wire [18:0] VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1;
VMStubs #("Tracklet") VMS_L5D3PHI2X2n4(
.data_in(VMR_L5D3_VMS_L5D3PHI2X2n4),
.enable(VMR_L5D3_VMS_L5D3PHI2X2n4_wr_en),
.number_out(VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1_number),
.read_add(VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1_read_add),
.data_out(VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X1n1;
wire VMR_L6D4_VMS_L6D4PHI3X1n1_wr_en;
wire [5:0] VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1_number;
wire [10:0] VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1_read_add;
wire [18:0] VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1;
VMStubs #("Tracklet") VMS_L6D4PHI3X1n1(
.data_in(VMR_L6D4_VMS_L6D4PHI3X1n1),
.enable(VMR_L6D4_VMS_L6D4PHI3X1n1_wr_en),
.number_out(VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1_number),
.read_add(VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1_read_add),
.data_out(VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X2n3;
wire VMR_L5D3_VMS_L5D3PHI3X2n3_wr_en;
wire [5:0] VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1_number;
wire [10:0] VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1_read_add;
wire [18:0] VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1;
VMStubs #("Tracklet") VMS_L5D3PHI3X2n3(
.data_in(VMR_L5D3_VMS_L5D3PHI3X2n3),
.enable(VMR_L5D3_VMS_L5D3PHI3X2n3_wr_en),
.number_out(VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1_number),
.read_add(VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1_read_add),
.data_out(VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X1n2;
wire VMR_L6D4_VMS_L6D4PHI3X1n2_wr_en;
wire [5:0] VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1_number;
wire [10:0] VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1_read_add;
wire [18:0] VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1;
VMStubs #("Tracklet") VMS_L6D4PHI3X1n2(
.data_in(VMR_L6D4_VMS_L6D4PHI3X1n2),
.enable(VMR_L6D4_VMS_L6D4PHI3X1n2_wr_en),
.number_out(VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1_number),
.read_add(VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1_read_add),
.data_out(VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X2n4;
wire VMR_L5D3_VMS_L5D3PHI3X2n4_wr_en;
wire [5:0] VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1_number;
wire [10:0] VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1_read_add;
wire [18:0] VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1;
VMStubs #("Tracklet") VMS_L5D3PHI3X2n4(
.data_in(VMR_L5D3_VMS_L5D3PHI3X2n4),
.enable(VMR_L5D3_VMS_L5D3PHI3X2n4_wr_en),
.number_out(VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1_number),
.read_add(VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1_read_add),
.data_out(VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI4X1n1;
wire VMR_L6D4_VMS_L6D4PHI4X1n1_wr_en;
wire [5:0] VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1_number;
wire [10:0] VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1_read_add;
wire [18:0] VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1;
VMStubs #("Tracklet") VMS_L6D4PHI4X1n1(
.data_in(VMR_L6D4_VMS_L6D4PHI4X1n1),
.enable(VMR_L6D4_VMS_L6D4PHI4X1n1_wr_en),
.number_out(VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1_number),
.read_add(VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1_read_add),
.data_out(VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI4X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X1n1;
wire VMR_L5D4_VMS_L5D4PHI1X1n1_wr_en;
wire [5:0] VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1_number;
wire [10:0] VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1_read_add;
wire [18:0] VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1;
VMStubs #("Tracklet") VMS_L5D4PHI1X1n1(
.data_in(VMR_L5D4_VMS_L5D4PHI1X1n1),
.enable(VMR_L5D4_VMS_L5D4PHI1X1n1_wr_en),
.number_out(VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1_number),
.read_add(VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1_read_add),
.data_out(VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI1X1n2;
wire VMR_L6D4_VMS_L6D4PHI1X1n2_wr_en;
wire [5:0] VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1_number;
wire [10:0] VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1_read_add;
wire [18:0] VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1;
VMStubs #("Tracklet") VMS_L6D4PHI1X1n2(
.data_in(VMR_L6D4_VMS_L6D4PHI1X1n2),
.enable(VMR_L6D4_VMS_L6D4PHI1X1n2_wr_en),
.number_out(VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1_number),
.read_add(VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1_read_add),
.data_out(VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X1n2;
wire VMR_L5D4_VMS_L5D4PHI1X1n2_wr_en;
wire [5:0] VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1_number;
wire [10:0] VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1_read_add;
wire [18:0] VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1;
VMStubs #("Tracklet") VMS_L5D4PHI1X1n2(
.data_in(VMR_L5D4_VMS_L5D4PHI1X1n2),
.enable(VMR_L5D4_VMS_L5D4PHI1X1n2_wr_en),
.number_out(VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1_number),
.read_add(VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1_read_add),
.data_out(VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X1n3;
wire VMR_L6D4_VMS_L6D4PHI2X1n3_wr_en;
wire [5:0] VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1_number;
wire [10:0] VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1_read_add;
wire [18:0] VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1;
VMStubs #("Tracklet") VMS_L6D4PHI2X1n3(
.data_in(VMR_L6D4_VMS_L6D4PHI2X1n3),
.enable(VMR_L6D4_VMS_L6D4PHI2X1n3_wr_en),
.number_out(VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1_number),
.read_add(VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1_read_add),
.data_out(VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X1n1;
wire VMR_L5D4_VMS_L5D4PHI2X1n1_wr_en;
wire [5:0] VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1_number;
wire [10:0] VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1_read_add;
wire [18:0] VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1;
VMStubs #("Tracklet") VMS_L5D4PHI2X1n1(
.data_in(VMR_L5D4_VMS_L5D4PHI2X1n1),
.enable(VMR_L5D4_VMS_L5D4PHI2X1n1_wr_en),
.number_out(VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1_number),
.read_add(VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1_read_add),
.data_out(VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X1n4;
wire VMR_L6D4_VMS_L6D4PHI2X1n4_wr_en;
wire [5:0] VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1_number;
wire [10:0] VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1_read_add;
wire [18:0] VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1;
VMStubs #("Tracklet") VMS_L6D4PHI2X1n4(
.data_in(VMR_L6D4_VMS_L6D4PHI2X1n4),
.enable(VMR_L6D4_VMS_L6D4PHI2X1n4_wr_en),
.number_out(VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1_number),
.read_add(VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1_read_add),
.data_out(VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X1n2;
wire VMR_L5D4_VMS_L5D4PHI2X1n2_wr_en;
wire [5:0] VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1_number;
wire [10:0] VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1_read_add;
wire [18:0] VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1;
VMStubs #("Tracklet") VMS_L5D4PHI2X1n2(
.data_in(VMR_L5D4_VMS_L5D4PHI2X1n2),
.enable(VMR_L5D4_VMS_L5D4PHI2X1n2_wr_en),
.number_out(VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1_number),
.read_add(VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1_read_add),
.data_out(VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X1n3;
wire VMR_L6D4_VMS_L6D4PHI3X1n3_wr_en;
wire [5:0] VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1_number;
wire [10:0] VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1_read_add;
wire [18:0] VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1;
VMStubs #("Tracklet") VMS_L6D4PHI3X1n3(
.data_in(VMR_L6D4_VMS_L6D4PHI3X1n3),
.enable(VMR_L6D4_VMS_L6D4PHI3X1n3_wr_en),
.number_out(VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1_number),
.read_add(VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1_read_add),
.data_out(VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X1n1;
wire VMR_L5D4_VMS_L5D4PHI3X1n1_wr_en;
wire [5:0] VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1_number;
wire [10:0] VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1_read_add;
wire [18:0] VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1;
VMStubs #("Tracklet") VMS_L5D4PHI3X1n1(
.data_in(VMR_L5D4_VMS_L5D4PHI3X1n1),
.enable(VMR_L5D4_VMS_L5D4PHI3X1n1_wr_en),
.number_out(VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1_number),
.read_add(VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1_read_add),
.data_out(VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X1n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X1n4;
wire VMR_L6D4_VMS_L6D4PHI3X1n4_wr_en;
wire [5:0] VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1_number;
wire [10:0] VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1_read_add;
wire [18:0] VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1;
VMStubs #("Tracklet") VMS_L6D4PHI3X1n4(
.data_in(VMR_L6D4_VMS_L6D4PHI3X1n4),
.enable(VMR_L6D4_VMS_L6D4PHI3X1n4_wr_en),
.number_out(VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1_number),
.read_add(VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1_read_add),
.data_out(VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X1n2;
wire VMR_L5D4_VMS_L5D4PHI3X1n2_wr_en;
wire [5:0] VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_number;
wire [10:0] VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_read_add;
wire [18:0] VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1;
VMStubs #("Tracklet") VMS_L5D4PHI3X1n2(
.data_in(VMR_L5D4_VMS_L5D4PHI3X1n2),
.enable(VMR_L5D4_VMS_L5D4PHI3X1n2_wr_en),
.number_out(VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_number),
.read_add(VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_read_add),
.data_out(VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI4X1n2;
wire VMR_L6D4_VMS_L6D4PHI4X1n2_wr_en;
wire [5:0] VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_number;
wire [10:0] VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_read_add;
wire [18:0] VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1;
VMStubs #("Tracklet") VMS_L6D4PHI4X1n2(
.data_in(VMR_L6D4_VMS_L6D4PHI4X1n2),
.enable(VMR_L6D4_VMS_L6D4PHI4X1n2_wr_en),
.number_out(VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_number),
.read_add(VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_read_add),
.data_out(VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X1n3;
wire VMR_L5D4_VMS_L5D4PHI1X1n3_wr_en;
wire [5:0] VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2_number;
wire [10:0] VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2_read_add;
wire [18:0] VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2;
VMStubs #("Tracklet") VMS_L5D4PHI1X1n3(
.data_in(VMR_L5D4_VMS_L5D4PHI1X1n3),
.enable(VMR_L5D4_VMS_L5D4PHI1X1n3_wr_en),
.number_out(VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2_number),
.read_add(VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2_read_add),
.data_out(VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI1X2n1;
wire VMR_L6D4_VMS_L6D4PHI1X2n1_wr_en;
wire [5:0] VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2_number;
wire [10:0] VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2_read_add;
wire [18:0] VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2;
VMStubs #("Tracklet") VMS_L6D4PHI1X2n1(
.data_in(VMR_L6D4_VMS_L6D4PHI1X2n1),
.enable(VMR_L6D4_VMS_L6D4PHI1X2n1_wr_en),
.number_out(VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2_number),
.read_add(VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2_read_add),
.data_out(VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X1n4;
wire VMR_L5D4_VMS_L5D4PHI1X1n4_wr_en;
wire [5:0] VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2_number;
wire [10:0] VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2_read_add;
wire [18:0] VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2;
VMStubs #("Tracklet") VMS_L5D4PHI1X1n4(
.data_in(VMR_L5D4_VMS_L5D4PHI1X1n4),
.enable(VMR_L5D4_VMS_L5D4PHI1X1n4_wr_en),
.number_out(VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2_number),
.read_add(VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2_read_add),
.data_out(VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X2n1;
wire VMR_L6D4_VMS_L6D4PHI2X2n1_wr_en;
wire [5:0] VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2_number;
wire [10:0] VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2_read_add;
wire [18:0] VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2;
VMStubs #("Tracklet") VMS_L6D4PHI2X2n1(
.data_in(VMR_L6D4_VMS_L6D4PHI2X2n1),
.enable(VMR_L6D4_VMS_L6D4PHI2X2n1_wr_en),
.number_out(VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2_number),
.read_add(VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2_read_add),
.data_out(VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X1n3;
wire VMR_L5D4_VMS_L5D4PHI2X1n3_wr_en;
wire [5:0] VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2_number;
wire [10:0] VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2_read_add;
wire [18:0] VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2;
VMStubs #("Tracklet") VMS_L5D4PHI2X1n3(
.data_in(VMR_L5D4_VMS_L5D4PHI2X1n3),
.enable(VMR_L5D4_VMS_L5D4PHI2X1n3_wr_en),
.number_out(VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2_number),
.read_add(VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2_read_add),
.data_out(VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X2n2;
wire VMR_L6D4_VMS_L6D4PHI2X2n2_wr_en;
wire [5:0] VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2_number;
wire [10:0] VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2_read_add;
wire [18:0] VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2;
VMStubs #("Tracklet") VMS_L6D4PHI2X2n2(
.data_in(VMR_L6D4_VMS_L6D4PHI2X2n2),
.enable(VMR_L6D4_VMS_L6D4PHI2X2n2_wr_en),
.number_out(VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2_number),
.read_add(VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2_read_add),
.data_out(VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X1n4;
wire VMR_L5D4_VMS_L5D4PHI2X1n4_wr_en;
wire [5:0] VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2_number;
wire [10:0] VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2_read_add;
wire [18:0] VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2;
VMStubs #("Tracklet") VMS_L5D4PHI2X1n4(
.data_in(VMR_L5D4_VMS_L5D4PHI2X1n4),
.enable(VMR_L5D4_VMS_L5D4PHI2X1n4_wr_en),
.number_out(VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2_number),
.read_add(VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2_read_add),
.data_out(VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X2n1;
wire VMR_L6D4_VMS_L6D4PHI3X2n1_wr_en;
wire [5:0] VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2_number;
wire [10:0] VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2_read_add;
wire [18:0] VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2;
VMStubs #("Tracklet") VMS_L6D4PHI3X2n1(
.data_in(VMR_L6D4_VMS_L6D4PHI3X2n1),
.enable(VMR_L6D4_VMS_L6D4PHI3X2n1_wr_en),
.number_out(VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2_number),
.read_add(VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2_read_add),
.data_out(VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X1n3;
wire VMR_L5D4_VMS_L5D4PHI3X1n3_wr_en;
wire [5:0] VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2_number;
wire [10:0] VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2_read_add;
wire [18:0] VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2;
VMStubs #("Tracklet") VMS_L5D4PHI3X1n3(
.data_in(VMR_L5D4_VMS_L5D4PHI3X1n3),
.enable(VMR_L5D4_VMS_L5D4PHI3X1n3_wr_en),
.number_out(VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2_number),
.read_add(VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2_read_add),
.data_out(VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X2n2;
wire VMR_L6D4_VMS_L6D4PHI3X2n2_wr_en;
wire [5:0] VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2_number;
wire [10:0] VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2_read_add;
wire [18:0] VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2;
VMStubs #("Tracklet") VMS_L6D4PHI3X2n2(
.data_in(VMR_L6D4_VMS_L6D4PHI3X2n2),
.enable(VMR_L6D4_VMS_L6D4PHI3X2n2_wr_en),
.number_out(VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2_number),
.read_add(VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2_read_add),
.data_out(VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X1n4;
wire VMR_L5D4_VMS_L5D4PHI3X1n4_wr_en;
wire [5:0] VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2_number;
wire [10:0] VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2_read_add;
wire [18:0] VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2;
VMStubs #("Tracklet") VMS_L5D4PHI3X1n4(
.data_in(VMR_L5D4_VMS_L5D4PHI3X1n4),
.enable(VMR_L5D4_VMS_L5D4PHI3X1n4_wr_en),
.number_out(VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2_number),
.read_add(VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2_read_add),
.data_out(VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI4X2n1;
wire VMR_L6D4_VMS_L6D4PHI4X2n1_wr_en;
wire [5:0] VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2_number;
wire [10:0] VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2_read_add;
wire [18:0] VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2;
VMStubs #("Tracklet") VMS_L6D4PHI4X2n1(
.data_in(VMR_L6D4_VMS_L6D4PHI4X2n1),
.enable(VMR_L6D4_VMS_L6D4PHI4X2n1_wr_en),
.number_out(VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2_number),
.read_add(VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2_read_add),
.data_out(VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI4X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X2n1;
wire VMR_L5D4_VMS_L5D4PHI1X2n1_wr_en;
wire [5:0] VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2_number;
wire [10:0] VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2_read_add;
wire [18:0] VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2;
VMStubs #("Tracklet") VMS_L5D4PHI1X2n1(
.data_in(VMR_L5D4_VMS_L5D4PHI1X2n1),
.enable(VMR_L5D4_VMS_L5D4PHI1X2n1_wr_en),
.number_out(VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2_number),
.read_add(VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2_read_add),
.data_out(VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI1X2n2;
wire VMR_L6D4_VMS_L6D4PHI1X2n2_wr_en;
wire [5:0] VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2_number;
wire [10:0] VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2_read_add;
wire [18:0] VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2;
VMStubs #("Tracklet") VMS_L6D4PHI1X2n2(
.data_in(VMR_L6D4_VMS_L6D4PHI1X2n2),
.enable(VMR_L6D4_VMS_L6D4PHI1X2n2_wr_en),
.number_out(VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2_number),
.read_add(VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2_read_add),
.data_out(VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X2n2;
wire VMR_L5D4_VMS_L5D4PHI1X2n2_wr_en;
wire [5:0] VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2_number;
wire [10:0] VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2_read_add;
wire [18:0] VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2;
VMStubs #("Tracklet") VMS_L5D4PHI1X2n2(
.data_in(VMR_L5D4_VMS_L5D4PHI1X2n2),
.enable(VMR_L5D4_VMS_L5D4PHI1X2n2_wr_en),
.number_out(VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2_number),
.read_add(VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2_read_add),
.data_out(VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X2n3;
wire VMR_L6D4_VMS_L6D4PHI2X2n3_wr_en;
wire [5:0] VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2_number;
wire [10:0] VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2_read_add;
wire [18:0] VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2;
VMStubs #("Tracklet") VMS_L6D4PHI2X2n3(
.data_in(VMR_L6D4_VMS_L6D4PHI2X2n3),
.enable(VMR_L6D4_VMS_L6D4PHI2X2n3_wr_en),
.number_out(VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2_number),
.read_add(VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2_read_add),
.data_out(VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X2n1;
wire VMR_L5D4_VMS_L5D4PHI2X2n1_wr_en;
wire [5:0] VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2_number;
wire [10:0] VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2_read_add;
wire [18:0] VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2;
VMStubs #("Tracklet") VMS_L5D4PHI2X2n1(
.data_in(VMR_L5D4_VMS_L5D4PHI2X2n1),
.enable(VMR_L5D4_VMS_L5D4PHI2X2n1_wr_en),
.number_out(VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2_number),
.read_add(VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2_read_add),
.data_out(VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X2n4;
wire VMR_L6D4_VMS_L6D4PHI2X2n4_wr_en;
wire [5:0] VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2_number;
wire [10:0] VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2_read_add;
wire [18:0] VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2;
VMStubs #("Tracklet") VMS_L6D4PHI2X2n4(
.data_in(VMR_L6D4_VMS_L6D4PHI2X2n4),
.enable(VMR_L6D4_VMS_L6D4PHI2X2n4_wr_en),
.number_out(VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2_number),
.read_add(VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2_read_add),
.data_out(VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X2n2;
wire VMR_L5D4_VMS_L5D4PHI2X2n2_wr_en;
wire [5:0] VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2_number;
wire [10:0] VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2_read_add;
wire [18:0] VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2;
VMStubs #("Tracklet") VMS_L5D4PHI2X2n2(
.data_in(VMR_L5D4_VMS_L5D4PHI2X2n2),
.enable(VMR_L5D4_VMS_L5D4PHI2X2n2_wr_en),
.number_out(VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2_number),
.read_add(VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2_read_add),
.data_out(VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X2n3;
wire VMR_L6D4_VMS_L6D4PHI3X2n3_wr_en;
wire [5:0] VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2_number;
wire [10:0] VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2_read_add;
wire [18:0] VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2;
VMStubs #("Tracklet") VMS_L6D4PHI3X2n3(
.data_in(VMR_L6D4_VMS_L6D4PHI3X2n3),
.enable(VMR_L6D4_VMS_L6D4PHI3X2n3_wr_en),
.number_out(VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2_number),
.read_add(VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2_read_add),
.data_out(VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X2n1;
wire VMR_L5D4_VMS_L5D4PHI3X2n1_wr_en;
wire [5:0] VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2_number;
wire [10:0] VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2_read_add;
wire [18:0] VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2;
VMStubs #("Tracklet") VMS_L5D4PHI3X2n1(
.data_in(VMR_L5D4_VMS_L5D4PHI3X2n1),
.enable(VMR_L5D4_VMS_L5D4PHI3X2n1_wr_en),
.number_out(VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2_number),
.read_add(VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2_read_add),
.data_out(VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X2n4;
wire VMR_L6D4_VMS_L6D4PHI3X2n4_wr_en;
wire [5:0] VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2_number;
wire [10:0] VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2_read_add;
wire [18:0] VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2;
VMStubs #("Tracklet") VMS_L6D4PHI3X2n4(
.data_in(VMR_L6D4_VMS_L6D4PHI3X2n4),
.enable(VMR_L6D4_VMS_L6D4PHI3X2n4_wr_en),
.number_out(VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2_number),
.read_add(VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2_read_add),
.data_out(VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X2n2;
wire VMR_L5D4_VMS_L5D4PHI3X2n2_wr_en;
wire [5:0] VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_number;
wire [10:0] VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_read_add;
wire [18:0] VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2;
VMStubs #("Tracklet") VMS_L5D4PHI3X2n2(
.data_in(VMR_L5D4_VMS_L5D4PHI3X2n2),
.enable(VMR_L5D4_VMS_L5D4PHI3X2n2_wr_en),
.number_out(VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_number),
.read_add(VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_read_add),
.data_out(VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI4X2n2;
wire VMR_L6D4_VMS_L6D4PHI4X2n2_wr_en;
wire [5:0] VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_number;
wire [10:0] VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_read_add;
wire [18:0] VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2;
VMStubs #("Tracklet") VMS_L6D4PHI4X2n2(
.data_in(VMR_L6D4_VMS_L6D4PHI4X2n2),
.enable(VMR_L6D4_VMS_L6D4PHI4X2n2_wr_en),
.number_out(VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_number),
.read_add(VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_read_add),
.data_out(VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI4X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X1_L2D3PHI1X1_SP_L1D3PHI1X1_L2D3PHI1X1;
wire TE_L1D3PHI1X1_L2D3PHI1X1_SP_L1D3PHI1X1_L2D3PHI1X1_wr_en;
wire [5:0] SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1X1_L2D3PHI1X1(
.data_in(TE_L1D3PHI1X1_L2D3PHI1X1_SP_L1D3PHI1X1_L2D3PHI1X1),
.enable(TE_L1D3PHI1X1_L2D3PHI1X1_SP_L1D3PHI1X1_L2D3PHI1X1_wr_en),
.number_out(SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3),
.start(TE_L1D3PHI1X1_L2D3PHI1X1_start),
.done(SP_L1D3PHI1X1_L2D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X1_L2D3PHI2X1_SP_L1D3PHI1X1_L2D3PHI2X1;
wire TE_L1D3PHI1X1_L2D3PHI2X1_SP_L1D3PHI1X1_L2D3PHI2X1_wr_en;
wire [5:0] SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1X1_L2D3PHI2X1(
.data_in(TE_L1D3PHI1X1_L2D3PHI2X1_SP_L1D3PHI1X1_L2D3PHI2X1),
.enable(TE_L1D3PHI1X1_L2D3PHI2X1_SP_L1D3PHI1X1_L2D3PHI2X1_wr_en),
.number_out(SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3),
.start(TE_L1D3PHI1X1_L2D3PHI2X1_start),
.done(SP_L1D3PHI1X1_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X1_L2D3PHI2X1_SP_L1D3PHI2X1_L2D3PHI2X1;
wire TE_L1D3PHI2X1_L2D3PHI2X1_SP_L1D3PHI2X1_L2D3PHI2X1_wr_en;
wire [5:0] SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2X1_L2D3PHI2X1(
.data_in(TE_L1D3PHI2X1_L2D3PHI2X1_SP_L1D3PHI2X1_L2D3PHI2X1),
.enable(TE_L1D3PHI2X1_L2D3PHI2X1_SP_L1D3PHI2X1_L2D3PHI2X1_wr_en),
.number_out(SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3),
.start(TE_L1D3PHI2X1_L2D3PHI2X1_start),
.done(SP_L1D3PHI2X1_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X1_L2D3PHI3X1_SP_L1D3PHI2X1_L2D3PHI3X1;
wire TE_L1D3PHI2X1_L2D3PHI3X1_SP_L1D3PHI2X1_L2D3PHI3X1_wr_en;
wire [5:0] SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2X1_L2D3PHI3X1(
.data_in(TE_L1D3PHI2X1_L2D3PHI3X1_SP_L1D3PHI2X1_L2D3PHI3X1),
.enable(TE_L1D3PHI2X1_L2D3PHI3X1_SP_L1D3PHI2X1_L2D3PHI3X1_wr_en),
.number_out(SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3),
.start(TE_L1D3PHI2X1_L2D3PHI3X1_start),
.done(SP_L1D3PHI2X1_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X1_L2D3PHI3X1_SP_L1D3PHI3X1_L2D3PHI3X1;
wire TE_L1D3PHI3X1_L2D3PHI3X1_SP_L1D3PHI3X1_L2D3PHI3X1_wr_en;
wire [5:0] SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3X1_L2D3PHI3X1(
.data_in(TE_L1D3PHI3X1_L2D3PHI3X1_SP_L1D3PHI3X1_L2D3PHI3X1),
.enable(TE_L1D3PHI3X1_L2D3PHI3X1_SP_L1D3PHI3X1_L2D3PHI3X1_wr_en),
.number_out(SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3),
.start(TE_L1D3PHI3X1_L2D3PHI3X1_start),
.done(SP_L1D3PHI3X1_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X1_L2D3PHI4X1_SP_L1D3PHI3X1_L2D3PHI4X1;
wire TE_L1D3PHI3X1_L2D3PHI4X1_SP_L1D3PHI3X1_L2D3PHI4X1_wr_en;
wire [5:0] SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3X1_L2D3PHI4X1(
.data_in(TE_L1D3PHI3X1_L2D3PHI4X1_SP_L1D3PHI3X1_L2D3PHI4X1),
.enable(TE_L1D3PHI3X1_L2D3PHI4X1_SP_L1D3PHI3X1_L2D3PHI4X1_wr_en),
.number_out(SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3),
.start(TE_L1D3PHI3X1_L2D3PHI4X1_start),
.done(SP_L1D3PHI3X1_L2D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X1_L2D3PHI1X2_SP_L1D3PHI1X1_L2D3PHI1X2;
wire TE_L1D3PHI1X1_L2D3PHI1X2_SP_L1D3PHI1X1_L2D3PHI1X2_wr_en;
wire [5:0] SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1X1_L2D3PHI1X2(
.data_in(TE_L1D3PHI1X1_L2D3PHI1X2_SP_L1D3PHI1X1_L2D3PHI1X2),
.enable(TE_L1D3PHI1X1_L2D3PHI1X2_SP_L1D3PHI1X1_L2D3PHI1X2_wr_en),
.number_out(SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3),
.start(TE_L1D3PHI1X1_L2D3PHI1X2_start),
.done(SP_L1D3PHI1X1_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X1_L2D3PHI2X2_SP_L1D3PHI1X1_L2D3PHI2X2;
wire TE_L1D3PHI1X1_L2D3PHI2X2_SP_L1D3PHI1X1_L2D3PHI2X2_wr_en;
wire [5:0] SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1X1_L2D3PHI2X2(
.data_in(TE_L1D3PHI1X1_L2D3PHI2X2_SP_L1D3PHI1X1_L2D3PHI2X2),
.enable(TE_L1D3PHI1X1_L2D3PHI2X2_SP_L1D3PHI1X1_L2D3PHI2X2_wr_en),
.number_out(SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3),
.start(TE_L1D3PHI1X1_L2D3PHI2X2_start),
.done(SP_L1D3PHI1X1_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X1_L2D3PHI2X2_SP_L1D3PHI2X1_L2D3PHI2X2;
wire TE_L1D3PHI2X1_L2D3PHI2X2_SP_L1D3PHI2X1_L2D3PHI2X2_wr_en;
wire [5:0] SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2X1_L2D3PHI2X2(
.data_in(TE_L1D3PHI2X1_L2D3PHI2X2_SP_L1D3PHI2X1_L2D3PHI2X2),
.enable(TE_L1D3PHI2X1_L2D3PHI2X2_SP_L1D3PHI2X1_L2D3PHI2X2_wr_en),
.number_out(SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3),
.start(TE_L1D3PHI2X1_L2D3PHI2X2_start),
.done(SP_L1D3PHI2X1_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X1_L2D3PHI3X2_SP_L1D3PHI2X1_L2D3PHI3X2;
wire TE_L1D3PHI2X1_L2D3PHI3X2_SP_L1D3PHI2X1_L2D3PHI3X2_wr_en;
wire [5:0] SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2X1_L2D3PHI3X2(
.data_in(TE_L1D3PHI2X1_L2D3PHI3X2_SP_L1D3PHI2X1_L2D3PHI3X2),
.enable(TE_L1D3PHI2X1_L2D3PHI3X2_SP_L1D3PHI2X1_L2D3PHI3X2_wr_en),
.number_out(SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3),
.start(TE_L1D3PHI2X1_L2D3PHI3X2_start),
.done(SP_L1D3PHI2X1_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X1_L2D3PHI3X2_SP_L1D3PHI3X1_L2D3PHI3X2;
wire TE_L1D3PHI3X1_L2D3PHI3X2_SP_L1D3PHI3X1_L2D3PHI3X2_wr_en;
wire [5:0] SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3X1_L2D3PHI3X2(
.data_in(TE_L1D3PHI3X1_L2D3PHI3X2_SP_L1D3PHI3X1_L2D3PHI3X2),
.enable(TE_L1D3PHI3X1_L2D3PHI3X2_SP_L1D3PHI3X1_L2D3PHI3X2_wr_en),
.number_out(SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3),
.start(TE_L1D3PHI3X1_L2D3PHI3X2_start),
.done(SP_L1D3PHI3X1_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X1_L2D3PHI4X2_SP_L1D3PHI3X1_L2D3PHI4X2;
wire TE_L1D3PHI3X1_L2D3PHI4X2_SP_L1D3PHI3X1_L2D3PHI4X2_wr_en;
wire [5:0] SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3X1_L2D3PHI4X2(
.data_in(TE_L1D3PHI3X1_L2D3PHI4X2_SP_L1D3PHI3X1_L2D3PHI4X2),
.enable(TE_L1D3PHI3X1_L2D3PHI4X2_SP_L1D3PHI3X1_L2D3PHI4X2_wr_en),
.number_out(SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3),
.start(TE_L1D3PHI3X1_L2D3PHI4X2_start),
.done(SP_L1D3PHI3X1_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X2_L2D3PHI1X2_SP_L1D3PHI1X2_L2D3PHI1X2;
wire TE_L1D3PHI1X2_L2D3PHI1X2_SP_L1D3PHI1X2_L2D3PHI1X2_wr_en;
wire [5:0] SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1X2_L2D3PHI1X2(
.data_in(TE_L1D3PHI1X2_L2D3PHI1X2_SP_L1D3PHI1X2_L2D3PHI1X2),
.enable(TE_L1D3PHI1X2_L2D3PHI1X2_SP_L1D3PHI1X2_L2D3PHI1X2_wr_en),
.number_out(SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3),
.start(TE_L1D3PHI1X2_L2D3PHI1X2_start),
.done(SP_L1D3PHI1X2_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X2_L2D3PHI2X2_SP_L1D3PHI1X2_L2D3PHI2X2;
wire TE_L1D3PHI1X2_L2D3PHI2X2_SP_L1D3PHI1X2_L2D3PHI2X2_wr_en;
wire [5:0] SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI1X2_L2D3PHI2X2(
.data_in(TE_L1D3PHI1X2_L2D3PHI2X2_SP_L1D3PHI1X2_L2D3PHI2X2),
.enable(TE_L1D3PHI1X2_L2D3PHI2X2_SP_L1D3PHI1X2_L2D3PHI2X2_wr_en),
.number_out(SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3),
.start(TE_L1D3PHI1X2_L2D3PHI2X2_start),
.done(SP_L1D3PHI1X2_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X2_L2D3PHI2X2_SP_L1D3PHI2X2_L2D3PHI2X2;
wire TE_L1D3PHI2X2_L2D3PHI2X2_SP_L1D3PHI2X2_L2D3PHI2X2_wr_en;
wire [5:0] SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2X2_L2D3PHI2X2(
.data_in(TE_L1D3PHI2X2_L2D3PHI2X2_SP_L1D3PHI2X2_L2D3PHI2X2),
.enable(TE_L1D3PHI2X2_L2D3PHI2X2_SP_L1D3PHI2X2_L2D3PHI2X2_wr_en),
.number_out(SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3),
.start(TE_L1D3PHI2X2_L2D3PHI2X2_start),
.done(SP_L1D3PHI2X2_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X2_L2D3PHI3X2_SP_L1D3PHI2X2_L2D3PHI3X2;
wire TE_L1D3PHI2X2_L2D3PHI3X2_SP_L1D3PHI2X2_L2D3PHI3X2_wr_en;
wire [5:0] SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI2X2_L2D3PHI3X2(
.data_in(TE_L1D3PHI2X2_L2D3PHI3X2_SP_L1D3PHI2X2_L2D3PHI3X2),
.enable(TE_L1D3PHI2X2_L2D3PHI3X2_SP_L1D3PHI2X2_L2D3PHI3X2_wr_en),
.number_out(SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3),
.start(TE_L1D3PHI2X2_L2D3PHI3X2_start),
.done(SP_L1D3PHI2X2_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X2_L2D3PHI3X2_SP_L1D3PHI3X2_L2D3PHI3X2;
wire TE_L1D3PHI3X2_L2D3PHI3X2_SP_L1D3PHI3X2_L2D3PHI3X2_wr_en;
wire [5:0] SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3X2_L2D3PHI3X2(
.data_in(TE_L1D3PHI3X2_L2D3PHI3X2_SP_L1D3PHI3X2_L2D3PHI3X2),
.enable(TE_L1D3PHI3X2_L2D3PHI3X2_SP_L1D3PHI3X2_L2D3PHI3X2_wr_en),
.number_out(SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3),
.start(TE_L1D3PHI3X2_L2D3PHI3X2_start),
.done(SP_L1D3PHI3X2_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X2_L2D3PHI4X2_SP_L1D3PHI3X2_L2D3PHI4X2;
wire TE_L1D3PHI3X2_L2D3PHI4X2_SP_L1D3PHI3X2_L2D3PHI4X2_wr_en;
wire [5:0] SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3_number;
wire [8:0] SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3_read_add;
wire [11:0] SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3;
StubPairs  SP_L1D3PHI3X2_L2D3PHI4X2(
.data_in(TE_L1D3PHI3X2_L2D3PHI4X2_SP_L1D3PHI3X2_L2D3PHI4X2),
.enable(TE_L1D3PHI3X2_L2D3PHI4X2_SP_L1D3PHI3X2_L2D3PHI4X2_wr_en),
.number_out(SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3_number),
.read_add(SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3_read_add),
.data_out(SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3),
.start(TE_L1D3PHI3X2_L2D3PHI4X2_start),
.done(SP_L1D3PHI3X2_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L1D3_AS_L1D3n1;
wire VMR_L1D3_AS_L1D3n1_wr_en;
wire [10:0] AS_L1D3n1_TC_L1D3L2D3_read_add;
wire [35:0] AS_L1D3n1_TC_L1D3L2D3;
AllStubs  AS_L1D3n1(
.data_in(VMR_L1D3_AS_L1D3n1),
.enable(VMR_L1D3_AS_L1D3n1_wr_en),
.read_add(AS_L1D3n1_TC_L1D3L2D3_read_add),
.data_out(AS_L1D3n1_TC_L1D3L2D3),
.start(VMR_L1D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L2D3_AS_L2D3n1;
wire VMR_L2D3_AS_L2D3n1_wr_en;
wire [10:0] AS_L2D3n1_TC_L1D3L2D3_read_add;
wire [35:0] AS_L2D3n1_TC_L1D3L2D3;
AllStubs  AS_L2D3n1(
.data_in(VMR_L2D3_AS_L2D3n1),
.enable(VMR_L2D3_AS_L2D3n1_wr_en),
.read_add(AS_L2D3n1_TC_L1D3L2D3_read_add),
.data_out(AS_L2D3n1_TC_L1D3L2D3),
.start(VMR_L2D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X1_L2D4PHI1X1_SP_L1D3PHI1X1_L2D4PHI1X1;
wire TE_L1D3PHI1X1_L2D4PHI1X1_SP_L1D3PHI1X1_L2D4PHI1X1_wr_en;
wire [5:0] SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1X1_L2D4PHI1X1(
.data_in(TE_L1D3PHI1X1_L2D4PHI1X1_SP_L1D3PHI1X1_L2D4PHI1X1),
.enable(TE_L1D3PHI1X1_L2D4PHI1X1_SP_L1D3PHI1X1_L2D4PHI1X1_wr_en),
.number_out(SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4),
.start(TE_L1D3PHI1X1_L2D4PHI1X1_start),
.done(SP_L1D3PHI1X1_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X1_L2D4PHI2X1_SP_L1D3PHI1X1_L2D4PHI2X1;
wire TE_L1D3PHI1X1_L2D4PHI2X1_SP_L1D3PHI1X1_L2D4PHI2X1_wr_en;
wire [5:0] SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1X1_L2D4PHI2X1(
.data_in(TE_L1D3PHI1X1_L2D4PHI2X1_SP_L1D3PHI1X1_L2D4PHI2X1),
.enable(TE_L1D3PHI1X1_L2D4PHI2X1_SP_L1D3PHI1X1_L2D4PHI2X1_wr_en),
.number_out(SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4),
.start(TE_L1D3PHI1X1_L2D4PHI2X1_start),
.done(SP_L1D3PHI1X1_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X1_L2D4PHI2X1_SP_L1D3PHI2X1_L2D4PHI2X1;
wire TE_L1D3PHI2X1_L2D4PHI2X1_SP_L1D3PHI2X1_L2D4PHI2X1_wr_en;
wire [5:0] SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2X1_L2D4PHI2X1(
.data_in(TE_L1D3PHI2X1_L2D4PHI2X1_SP_L1D3PHI2X1_L2D4PHI2X1),
.enable(TE_L1D3PHI2X1_L2D4PHI2X1_SP_L1D3PHI2X1_L2D4PHI2X1_wr_en),
.number_out(SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4),
.start(TE_L1D3PHI2X1_L2D4PHI2X1_start),
.done(SP_L1D3PHI2X1_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X1_L2D4PHI3X1_SP_L1D3PHI2X1_L2D4PHI3X1;
wire TE_L1D3PHI2X1_L2D4PHI3X1_SP_L1D3PHI2X1_L2D4PHI3X1_wr_en;
wire [5:0] SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2X1_L2D4PHI3X1(
.data_in(TE_L1D3PHI2X1_L2D4PHI3X1_SP_L1D3PHI2X1_L2D4PHI3X1),
.enable(TE_L1D3PHI2X1_L2D4PHI3X1_SP_L1D3PHI2X1_L2D4PHI3X1_wr_en),
.number_out(SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4),
.start(TE_L1D3PHI2X1_L2D4PHI3X1_start),
.done(SP_L1D3PHI2X1_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X1_L2D4PHI3X1_SP_L1D3PHI3X1_L2D4PHI3X1;
wire TE_L1D3PHI3X1_L2D4PHI3X1_SP_L1D3PHI3X1_L2D4PHI3X1_wr_en;
wire [5:0] SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3X1_L2D4PHI3X1(
.data_in(TE_L1D3PHI3X1_L2D4PHI3X1_SP_L1D3PHI3X1_L2D4PHI3X1),
.enable(TE_L1D3PHI3X1_L2D4PHI3X1_SP_L1D3PHI3X1_L2D4PHI3X1_wr_en),
.number_out(SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4),
.start(TE_L1D3PHI3X1_L2D4PHI3X1_start),
.done(SP_L1D3PHI3X1_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X1_L2D4PHI4X1_SP_L1D3PHI3X1_L2D4PHI4X1;
wire TE_L1D3PHI3X1_L2D4PHI4X1_SP_L1D3PHI3X1_L2D4PHI4X1_wr_en;
wire [5:0] SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3X1_L2D4PHI4X1(
.data_in(TE_L1D3PHI3X1_L2D4PHI4X1_SP_L1D3PHI3X1_L2D4PHI4X1),
.enable(TE_L1D3PHI3X1_L2D4PHI4X1_SP_L1D3PHI3X1_L2D4PHI4X1_wr_en),
.number_out(SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4),
.start(TE_L1D3PHI3X1_L2D4PHI4X1_start),
.done(SP_L1D3PHI3X1_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X2_L2D4PHI1X1_SP_L1D3PHI1X2_L2D4PHI1X1;
wire TE_L1D3PHI1X2_L2D4PHI1X1_SP_L1D3PHI1X2_L2D4PHI1X1_wr_en;
wire [5:0] SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1X2_L2D4PHI1X1(
.data_in(TE_L1D3PHI1X2_L2D4PHI1X1_SP_L1D3PHI1X2_L2D4PHI1X1),
.enable(TE_L1D3PHI1X2_L2D4PHI1X1_SP_L1D3PHI1X2_L2D4PHI1X1_wr_en),
.number_out(SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4),
.start(TE_L1D3PHI1X2_L2D4PHI1X1_start),
.done(SP_L1D3PHI1X2_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X2_L2D4PHI2X1_SP_L1D3PHI1X2_L2D4PHI2X1;
wire TE_L1D3PHI1X2_L2D4PHI2X1_SP_L1D3PHI1X2_L2D4PHI2X1_wr_en;
wire [5:0] SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1X2_L2D4PHI2X1(
.data_in(TE_L1D3PHI1X2_L2D4PHI2X1_SP_L1D3PHI1X2_L2D4PHI2X1),
.enable(TE_L1D3PHI1X2_L2D4PHI2X1_SP_L1D3PHI1X2_L2D4PHI2X1_wr_en),
.number_out(SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4),
.start(TE_L1D3PHI1X2_L2D4PHI2X1_start),
.done(SP_L1D3PHI1X2_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X2_L2D4PHI2X1_SP_L1D3PHI2X2_L2D4PHI2X1;
wire TE_L1D3PHI2X2_L2D4PHI2X1_SP_L1D3PHI2X2_L2D4PHI2X1_wr_en;
wire [5:0] SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2X2_L2D4PHI2X1(
.data_in(TE_L1D3PHI2X2_L2D4PHI2X1_SP_L1D3PHI2X2_L2D4PHI2X1),
.enable(TE_L1D3PHI2X2_L2D4PHI2X1_SP_L1D3PHI2X2_L2D4PHI2X1_wr_en),
.number_out(SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4),
.start(TE_L1D3PHI2X2_L2D4PHI2X1_start),
.done(SP_L1D3PHI2X2_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X2_L2D4PHI3X1_SP_L1D3PHI2X2_L2D4PHI3X1;
wire TE_L1D3PHI2X2_L2D4PHI3X1_SP_L1D3PHI2X2_L2D4PHI3X1_wr_en;
wire [5:0] SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2X2_L2D4PHI3X1(
.data_in(TE_L1D3PHI2X2_L2D4PHI3X1_SP_L1D3PHI2X2_L2D4PHI3X1),
.enable(TE_L1D3PHI2X2_L2D4PHI3X1_SP_L1D3PHI2X2_L2D4PHI3X1_wr_en),
.number_out(SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4),
.start(TE_L1D3PHI2X2_L2D4PHI3X1_start),
.done(SP_L1D3PHI2X2_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X2_L2D4PHI3X1_SP_L1D3PHI3X2_L2D4PHI3X1;
wire TE_L1D3PHI3X2_L2D4PHI3X1_SP_L1D3PHI3X2_L2D4PHI3X1_wr_en;
wire [5:0] SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3X2_L2D4PHI3X1(
.data_in(TE_L1D3PHI3X2_L2D4PHI3X1_SP_L1D3PHI3X2_L2D4PHI3X1),
.enable(TE_L1D3PHI3X2_L2D4PHI3X1_SP_L1D3PHI3X2_L2D4PHI3X1_wr_en),
.number_out(SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4),
.start(TE_L1D3PHI3X2_L2D4PHI3X1_start),
.done(SP_L1D3PHI3X2_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X2_L2D4PHI4X1_SP_L1D3PHI3X2_L2D4PHI4X1;
wire TE_L1D3PHI3X2_L2D4PHI4X1_SP_L1D3PHI3X2_L2D4PHI4X1_wr_en;
wire [5:0] SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3X2_L2D4PHI4X1(
.data_in(TE_L1D3PHI3X2_L2D4PHI4X1_SP_L1D3PHI3X2_L2D4PHI4X1),
.enable(TE_L1D3PHI3X2_L2D4PHI4X1_SP_L1D3PHI3X2_L2D4PHI4X1_wr_en),
.number_out(SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4),
.start(TE_L1D3PHI3X2_L2D4PHI4X1_start),
.done(SP_L1D3PHI3X2_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X2_L2D4PHI1X2_SP_L1D3PHI1X2_L2D4PHI1X2;
wire TE_L1D3PHI1X2_L2D4PHI1X2_SP_L1D3PHI1X2_L2D4PHI1X2_wr_en;
wire [5:0] SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1X2_L2D4PHI1X2(
.data_in(TE_L1D3PHI1X2_L2D4PHI1X2_SP_L1D3PHI1X2_L2D4PHI1X2),
.enable(TE_L1D3PHI1X2_L2D4PHI1X2_SP_L1D3PHI1X2_L2D4PHI1X2_wr_en),
.number_out(SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4),
.start(TE_L1D3PHI1X2_L2D4PHI1X2_start),
.done(SP_L1D3PHI1X2_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI1X2_L2D4PHI2X2_SP_L1D3PHI1X2_L2D4PHI2X2;
wire TE_L1D3PHI1X2_L2D4PHI2X2_SP_L1D3PHI1X2_L2D4PHI2X2_wr_en;
wire [5:0] SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI1X2_L2D4PHI2X2(
.data_in(TE_L1D3PHI1X2_L2D4PHI2X2_SP_L1D3PHI1X2_L2D4PHI2X2),
.enable(TE_L1D3PHI1X2_L2D4PHI2X2_SP_L1D3PHI1X2_L2D4PHI2X2_wr_en),
.number_out(SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4),
.start(TE_L1D3PHI1X2_L2D4PHI2X2_start),
.done(SP_L1D3PHI1X2_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X2_L2D4PHI2X2_SP_L1D3PHI2X2_L2D4PHI2X2;
wire TE_L1D3PHI2X2_L2D4PHI2X2_SP_L1D3PHI2X2_L2D4PHI2X2_wr_en;
wire [5:0] SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2X2_L2D4PHI2X2(
.data_in(TE_L1D3PHI2X2_L2D4PHI2X2_SP_L1D3PHI2X2_L2D4PHI2X2),
.enable(TE_L1D3PHI2X2_L2D4PHI2X2_SP_L1D3PHI2X2_L2D4PHI2X2_wr_en),
.number_out(SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4),
.start(TE_L1D3PHI2X2_L2D4PHI2X2_start),
.done(SP_L1D3PHI2X2_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI2X2_L2D4PHI3X2_SP_L1D3PHI2X2_L2D4PHI3X2;
wire TE_L1D3PHI2X2_L2D4PHI3X2_SP_L1D3PHI2X2_L2D4PHI3X2_wr_en;
wire [5:0] SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI2X2_L2D4PHI3X2(
.data_in(TE_L1D3PHI2X2_L2D4PHI3X2_SP_L1D3PHI2X2_L2D4PHI3X2),
.enable(TE_L1D3PHI2X2_L2D4PHI3X2_SP_L1D3PHI2X2_L2D4PHI3X2_wr_en),
.number_out(SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4),
.start(TE_L1D3PHI2X2_L2D4PHI3X2_start),
.done(SP_L1D3PHI2X2_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X2_L2D4PHI3X2_SP_L1D3PHI3X2_L2D4PHI3X2;
wire TE_L1D3PHI3X2_L2D4PHI3X2_SP_L1D3PHI3X2_L2D4PHI3X2_wr_en;
wire [5:0] SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3X2_L2D4PHI3X2(
.data_in(TE_L1D3PHI3X2_L2D4PHI3X2_SP_L1D3PHI3X2_L2D4PHI3X2),
.enable(TE_L1D3PHI3X2_L2D4PHI3X2_SP_L1D3PHI3X2_L2D4PHI3X2_wr_en),
.number_out(SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4),
.start(TE_L1D3PHI3X2_L2D4PHI3X2_start),
.done(SP_L1D3PHI3X2_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D3PHI3X2_L2D4PHI4X2_SP_L1D3PHI3X2_L2D4PHI4X2;
wire TE_L1D3PHI3X2_L2D4PHI4X2_SP_L1D3PHI3X2_L2D4PHI4X2_wr_en;
wire [5:0] SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4_number;
wire [8:0] SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4_read_add;
wire [11:0] SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4;
StubPairs  SP_L1D3PHI3X2_L2D4PHI4X2(
.data_in(TE_L1D3PHI3X2_L2D4PHI4X2_SP_L1D3PHI3X2_L2D4PHI4X2),
.enable(TE_L1D3PHI3X2_L2D4PHI4X2_SP_L1D3PHI3X2_L2D4PHI4X2_wr_en),
.number_out(SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4_number),
.read_add(SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4_read_add),
.data_out(SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4),
.start(TE_L1D3PHI3X2_L2D4PHI4X2_start),
.done(SP_L1D3PHI3X2_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L1D3_AS_L1D3n2;
wire VMR_L1D3_AS_L1D3n2_wr_en;
wire [10:0] AS_L1D3n2_TC_L1D3L2D4_read_add;
wire [35:0] AS_L1D3n2_TC_L1D3L2D4;
AllStubs  AS_L1D3n2(
.data_in(VMR_L1D3_AS_L1D3n2),
.enable(VMR_L1D3_AS_L1D3n2_wr_en),
.read_add(AS_L1D3n2_TC_L1D3L2D4_read_add),
.data_out(AS_L1D3n2_TC_L1D3L2D4),
.start(VMR_L1D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L2D4_AS_L2D4n1;
wire VMR_L2D4_AS_L2D4n1_wr_en;
wire [10:0] AS_L2D4n1_TC_L1D3L2D4_read_add;
wire [35:0] AS_L2D4n1_TC_L1D3L2D4;
AllStubs  AS_L2D4n1(
.data_in(VMR_L2D4_AS_L2D4n1),
.enable(VMR_L2D4_AS_L2D4n1_wr_en),
.read_add(AS_L2D4n1_TC_L1D3L2D4_read_add),
.data_out(AS_L2D4n1_TC_L1D3L2D4),
.start(VMR_L2D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D4PHI1X1_L2D4PHI1X2_SP_L1D4PHI1X1_L2D4PHI1X2;
wire TE_L1D4PHI1X1_L2D4PHI1X2_SP_L1D4PHI1X1_L2D4PHI1X2_wr_en;
wire [5:0] SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI1X1_L2D4PHI1X2(
.data_in(TE_L1D4PHI1X1_L2D4PHI1X2_SP_L1D4PHI1X1_L2D4PHI1X2),
.enable(TE_L1D4PHI1X1_L2D4PHI1X2_SP_L1D4PHI1X1_L2D4PHI1X2_wr_en),
.number_out(SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4),
.start(TE_L1D4PHI1X1_L2D4PHI1X2_start),
.done(SP_L1D4PHI1X1_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D4PHI1X1_L2D4PHI2X2_SP_L1D4PHI1X1_L2D4PHI2X2;
wire TE_L1D4PHI1X1_L2D4PHI2X2_SP_L1D4PHI1X1_L2D4PHI2X2_wr_en;
wire [5:0] SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI1X1_L2D4PHI2X2(
.data_in(TE_L1D4PHI1X1_L2D4PHI2X2_SP_L1D4PHI1X1_L2D4PHI2X2),
.enable(TE_L1D4PHI1X1_L2D4PHI2X2_SP_L1D4PHI1X1_L2D4PHI2X2_wr_en),
.number_out(SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4),
.start(TE_L1D4PHI1X1_L2D4PHI2X2_start),
.done(SP_L1D4PHI1X1_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D4PHI2X1_L2D4PHI2X2_SP_L1D4PHI2X1_L2D4PHI2X2;
wire TE_L1D4PHI2X1_L2D4PHI2X2_SP_L1D4PHI2X1_L2D4PHI2X2_wr_en;
wire [5:0] SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI2X1_L2D4PHI2X2(
.data_in(TE_L1D4PHI2X1_L2D4PHI2X2_SP_L1D4PHI2X1_L2D4PHI2X2),
.enable(TE_L1D4PHI2X1_L2D4PHI2X2_SP_L1D4PHI2X1_L2D4PHI2X2_wr_en),
.number_out(SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4),
.start(TE_L1D4PHI2X1_L2D4PHI2X2_start),
.done(SP_L1D4PHI2X1_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D4PHI2X1_L2D4PHI3X2_SP_L1D4PHI2X1_L2D4PHI3X2;
wire TE_L1D4PHI2X1_L2D4PHI3X2_SP_L1D4PHI2X1_L2D4PHI3X2_wr_en;
wire [5:0] SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI2X1_L2D4PHI3X2(
.data_in(TE_L1D4PHI2X1_L2D4PHI3X2_SP_L1D4PHI2X1_L2D4PHI3X2),
.enable(TE_L1D4PHI2X1_L2D4PHI3X2_SP_L1D4PHI2X1_L2D4PHI3X2_wr_en),
.number_out(SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4),
.start(TE_L1D4PHI2X1_L2D4PHI3X2_start),
.done(SP_L1D4PHI2X1_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D4PHI3X1_L2D4PHI3X2_SP_L1D4PHI3X1_L2D4PHI3X2;
wire TE_L1D4PHI3X1_L2D4PHI3X2_SP_L1D4PHI3X1_L2D4PHI3X2_wr_en;
wire [5:0] SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI3X1_L2D4PHI3X2(
.data_in(TE_L1D4PHI3X1_L2D4PHI3X2_SP_L1D4PHI3X1_L2D4PHI3X2),
.enable(TE_L1D4PHI3X1_L2D4PHI3X2_SP_L1D4PHI3X1_L2D4PHI3X2_wr_en),
.number_out(SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4),
.start(TE_L1D4PHI3X1_L2D4PHI3X2_start),
.done(SP_L1D4PHI3X1_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L1D4PHI3X1_L2D4PHI4X2_SP_L1D4PHI3X1_L2D4PHI4X2;
wire TE_L1D4PHI3X1_L2D4PHI4X2_SP_L1D4PHI3X1_L2D4PHI4X2_wr_en;
wire [5:0] SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4_number;
wire [8:0] SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4_read_add;
wire [11:0] SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4;
StubPairs  SP_L1D4PHI3X1_L2D4PHI4X2(
.data_in(TE_L1D4PHI3X1_L2D4PHI4X2_SP_L1D4PHI3X1_L2D4PHI4X2),
.enable(TE_L1D4PHI3X1_L2D4PHI4X2_SP_L1D4PHI3X1_L2D4PHI4X2_wr_en),
.number_out(SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4_number),
.read_add(SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4_read_add),
.data_out(SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4),
.start(TE_L1D4PHI3X1_L2D4PHI4X2_start),
.done(SP_L1D4PHI3X1_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L1D4_AS_L1D4n1;
wire VMR_L1D4_AS_L1D4n1_wr_en;
wire [10:0] AS_L1D4n1_TC_L1D4L2D4_read_add;
wire [35:0] AS_L1D4n1_TC_L1D4L2D4;
AllStubs  AS_L1D4n1(
.data_in(VMR_L1D4_AS_L1D4n1),
.enable(VMR_L1D4_AS_L1D4n1_wr_en),
.read_add(AS_L1D4n1_TC_L1D4L2D4_read_add),
.data_out(AS_L1D4n1_TC_L1D4L2D4),
.start(VMR_L1D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L2D4_AS_L2D4n2;
wire VMR_L2D4_AS_L2D4n2_wr_en;
wire [10:0] AS_L2D4n2_TC_L1D4L2D4_read_add;
wire [35:0] AS_L2D4n2_TC_L1D4L2D4;
AllStubs  AS_L2D4n2(
.data_in(VMR_L2D4_AS_L2D4n2),
.enable(VMR_L2D4_AS_L2D4n2_wr_en),
.read_add(AS_L2D4n2_TC_L1D4L2D4_read_add),
.data_out(AS_L2D4n2_TC_L1D4L2D4),
.start(VMR_L2D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI1X1_L4D3PHI1X1_SP_L3D3PHI1X1_L4D3PHI1X1;
wire TE_L3D3PHI1X1_L4D3PHI1X1_SP_L3D3PHI1X1_L4D3PHI1X1_wr_en;
wire [5:0] SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1X1_L4D3PHI1X1(
.data_in(TE_L3D3PHI1X1_L4D3PHI1X1_SP_L3D3PHI1X1_L4D3PHI1X1),
.enable(TE_L3D3PHI1X1_L4D3PHI1X1_SP_L3D3PHI1X1_L4D3PHI1X1_wr_en),
.number_out(SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3),
.start(TE_L3D3PHI1X1_L4D3PHI1X1_start),
.done(SP_L3D3PHI1X1_L4D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI1X1_L4D3PHI2X1_SP_L3D3PHI1X1_L4D3PHI2X1;
wire TE_L3D3PHI1X1_L4D3PHI2X1_SP_L3D3PHI1X1_L4D3PHI2X1_wr_en;
wire [5:0] SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1X1_L4D3PHI2X1(
.data_in(TE_L3D3PHI1X1_L4D3PHI2X1_SP_L3D3PHI1X1_L4D3PHI2X1),
.enable(TE_L3D3PHI1X1_L4D3PHI2X1_SP_L3D3PHI1X1_L4D3PHI2X1_wr_en),
.number_out(SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3),
.start(TE_L3D3PHI1X1_L4D3PHI2X1_start),
.done(SP_L3D3PHI1X1_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI2X1_L4D3PHI2X1_SP_L3D3PHI2X1_L4D3PHI2X1;
wire TE_L3D3PHI2X1_L4D3PHI2X1_SP_L3D3PHI2X1_L4D3PHI2X1_wr_en;
wire [5:0] SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2X1_L4D3PHI2X1(
.data_in(TE_L3D3PHI2X1_L4D3PHI2X1_SP_L3D3PHI2X1_L4D3PHI2X1),
.enable(TE_L3D3PHI2X1_L4D3PHI2X1_SP_L3D3PHI2X1_L4D3PHI2X1_wr_en),
.number_out(SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3),
.start(TE_L3D3PHI2X1_L4D3PHI2X1_start),
.done(SP_L3D3PHI2X1_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI2X1_L4D3PHI3X1_SP_L3D3PHI2X1_L4D3PHI3X1;
wire TE_L3D3PHI2X1_L4D3PHI3X1_SP_L3D3PHI2X1_L4D3PHI3X1_wr_en;
wire [5:0] SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2X1_L4D3PHI3X1(
.data_in(TE_L3D3PHI2X1_L4D3PHI3X1_SP_L3D3PHI2X1_L4D3PHI3X1),
.enable(TE_L3D3PHI2X1_L4D3PHI3X1_SP_L3D3PHI2X1_L4D3PHI3X1_wr_en),
.number_out(SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3),
.start(TE_L3D3PHI2X1_L4D3PHI3X1_start),
.done(SP_L3D3PHI2X1_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI3X1_L4D3PHI3X1_SP_L3D3PHI3X1_L4D3PHI3X1;
wire TE_L3D3PHI3X1_L4D3PHI3X1_SP_L3D3PHI3X1_L4D3PHI3X1_wr_en;
wire [5:0] SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3X1_L4D3PHI3X1(
.data_in(TE_L3D3PHI3X1_L4D3PHI3X1_SP_L3D3PHI3X1_L4D3PHI3X1),
.enable(TE_L3D3PHI3X1_L4D3PHI3X1_SP_L3D3PHI3X1_L4D3PHI3X1_wr_en),
.number_out(SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3),
.start(TE_L3D3PHI3X1_L4D3PHI3X1_start),
.done(SP_L3D3PHI3X1_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI3X1_L4D3PHI4X1_SP_L3D3PHI3X1_L4D3PHI4X1;
wire TE_L3D3PHI3X1_L4D3PHI4X1_SP_L3D3PHI3X1_L4D3PHI4X1_wr_en;
wire [5:0] SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3X1_L4D3PHI4X1(
.data_in(TE_L3D3PHI3X1_L4D3PHI4X1_SP_L3D3PHI3X1_L4D3PHI4X1),
.enable(TE_L3D3PHI3X1_L4D3PHI4X1_SP_L3D3PHI3X1_L4D3PHI4X1_wr_en),
.number_out(SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3),
.start(TE_L3D3PHI3X1_L4D3PHI4X1_start),
.done(SP_L3D3PHI3X1_L4D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI1X1_L4D3PHI1X2_SP_L3D3PHI1X1_L4D3PHI1X2;
wire TE_L3D3PHI1X1_L4D3PHI1X2_SP_L3D3PHI1X1_L4D3PHI1X2_wr_en;
wire [5:0] SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1X1_L4D3PHI1X2(
.data_in(TE_L3D3PHI1X1_L4D3PHI1X2_SP_L3D3PHI1X1_L4D3PHI1X2),
.enable(TE_L3D3PHI1X1_L4D3PHI1X2_SP_L3D3PHI1X1_L4D3PHI1X2_wr_en),
.number_out(SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3),
.start(TE_L3D3PHI1X1_L4D3PHI1X2_start),
.done(SP_L3D3PHI1X1_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI1X1_L4D3PHI2X2_SP_L3D3PHI1X1_L4D3PHI2X2;
wire TE_L3D3PHI1X1_L4D3PHI2X2_SP_L3D3PHI1X1_L4D3PHI2X2_wr_en;
wire [5:0] SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1X1_L4D3PHI2X2(
.data_in(TE_L3D3PHI1X1_L4D3PHI2X2_SP_L3D3PHI1X1_L4D3PHI2X2),
.enable(TE_L3D3PHI1X1_L4D3PHI2X2_SP_L3D3PHI1X1_L4D3PHI2X2_wr_en),
.number_out(SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3),
.start(TE_L3D3PHI1X1_L4D3PHI2X2_start),
.done(SP_L3D3PHI1X1_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI2X1_L4D3PHI2X2_SP_L3D3PHI2X1_L4D3PHI2X2;
wire TE_L3D3PHI2X1_L4D3PHI2X2_SP_L3D3PHI2X1_L4D3PHI2X2_wr_en;
wire [5:0] SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2X1_L4D3PHI2X2(
.data_in(TE_L3D3PHI2X1_L4D3PHI2X2_SP_L3D3PHI2X1_L4D3PHI2X2),
.enable(TE_L3D3PHI2X1_L4D3PHI2X2_SP_L3D3PHI2X1_L4D3PHI2X2_wr_en),
.number_out(SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3),
.start(TE_L3D3PHI2X1_L4D3PHI2X2_start),
.done(SP_L3D3PHI2X1_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI2X1_L4D3PHI3X2_SP_L3D3PHI2X1_L4D3PHI3X2;
wire TE_L3D3PHI2X1_L4D3PHI3X2_SP_L3D3PHI2X1_L4D3PHI3X2_wr_en;
wire [5:0] SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2X1_L4D3PHI3X2(
.data_in(TE_L3D3PHI2X1_L4D3PHI3X2_SP_L3D3PHI2X1_L4D3PHI3X2),
.enable(TE_L3D3PHI2X1_L4D3PHI3X2_SP_L3D3PHI2X1_L4D3PHI3X2_wr_en),
.number_out(SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3),
.start(TE_L3D3PHI2X1_L4D3PHI3X2_start),
.done(SP_L3D3PHI2X1_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI3X1_L4D3PHI3X2_SP_L3D3PHI3X1_L4D3PHI3X2;
wire TE_L3D3PHI3X1_L4D3PHI3X2_SP_L3D3PHI3X1_L4D3PHI3X2_wr_en;
wire [5:0] SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3X1_L4D3PHI3X2(
.data_in(TE_L3D3PHI3X1_L4D3PHI3X2_SP_L3D3PHI3X1_L4D3PHI3X2),
.enable(TE_L3D3PHI3X1_L4D3PHI3X2_SP_L3D3PHI3X1_L4D3PHI3X2_wr_en),
.number_out(SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3),
.start(TE_L3D3PHI3X1_L4D3PHI3X2_start),
.done(SP_L3D3PHI3X1_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI3X1_L4D3PHI4X2_SP_L3D3PHI3X1_L4D3PHI4X2;
wire TE_L3D3PHI3X1_L4D3PHI4X2_SP_L3D3PHI3X1_L4D3PHI4X2_wr_en;
wire [5:0] SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3X1_L4D3PHI4X2(
.data_in(TE_L3D3PHI3X1_L4D3PHI4X2_SP_L3D3PHI3X1_L4D3PHI4X2),
.enable(TE_L3D3PHI3X1_L4D3PHI4X2_SP_L3D3PHI3X1_L4D3PHI4X2_wr_en),
.number_out(SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3),
.start(TE_L3D3PHI3X1_L4D3PHI4X2_start),
.done(SP_L3D3PHI3X1_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI1X2_L4D3PHI1X2_SP_L3D3PHI1X2_L4D3PHI1X2;
wire TE_L3D3PHI1X2_L4D3PHI1X2_SP_L3D3PHI1X2_L4D3PHI1X2_wr_en;
wire [5:0] SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1X2_L4D3PHI1X2(
.data_in(TE_L3D3PHI1X2_L4D3PHI1X2_SP_L3D3PHI1X2_L4D3PHI1X2),
.enable(TE_L3D3PHI1X2_L4D3PHI1X2_SP_L3D3PHI1X2_L4D3PHI1X2_wr_en),
.number_out(SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3),
.start(TE_L3D3PHI1X2_L4D3PHI1X2_start),
.done(SP_L3D3PHI1X2_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI1X2_L4D3PHI2X2_SP_L3D3PHI1X2_L4D3PHI2X2;
wire TE_L3D3PHI1X2_L4D3PHI2X2_SP_L3D3PHI1X2_L4D3PHI2X2_wr_en;
wire [5:0] SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI1X2_L4D3PHI2X2(
.data_in(TE_L3D3PHI1X2_L4D3PHI2X2_SP_L3D3PHI1X2_L4D3PHI2X2),
.enable(TE_L3D3PHI1X2_L4D3PHI2X2_SP_L3D3PHI1X2_L4D3PHI2X2_wr_en),
.number_out(SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3),
.start(TE_L3D3PHI1X2_L4D3PHI2X2_start),
.done(SP_L3D3PHI1X2_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI2X2_L4D3PHI2X2_SP_L3D3PHI2X2_L4D3PHI2X2;
wire TE_L3D3PHI2X2_L4D3PHI2X2_SP_L3D3PHI2X2_L4D3PHI2X2_wr_en;
wire [5:0] SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2X2_L4D3PHI2X2(
.data_in(TE_L3D3PHI2X2_L4D3PHI2X2_SP_L3D3PHI2X2_L4D3PHI2X2),
.enable(TE_L3D3PHI2X2_L4D3PHI2X2_SP_L3D3PHI2X2_L4D3PHI2X2_wr_en),
.number_out(SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3),
.start(TE_L3D3PHI2X2_L4D3PHI2X2_start),
.done(SP_L3D3PHI2X2_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI2X2_L4D3PHI3X2_SP_L3D3PHI2X2_L4D3PHI3X2;
wire TE_L3D3PHI2X2_L4D3PHI3X2_SP_L3D3PHI2X2_L4D3PHI3X2_wr_en;
wire [5:0] SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI2X2_L4D3PHI3X2(
.data_in(TE_L3D3PHI2X2_L4D3PHI3X2_SP_L3D3PHI2X2_L4D3PHI3X2),
.enable(TE_L3D3PHI2X2_L4D3PHI3X2_SP_L3D3PHI2X2_L4D3PHI3X2_wr_en),
.number_out(SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3),
.start(TE_L3D3PHI2X2_L4D3PHI3X2_start),
.done(SP_L3D3PHI2X2_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI3X2_L4D3PHI3X2_SP_L3D3PHI3X2_L4D3PHI3X2;
wire TE_L3D3PHI3X2_L4D3PHI3X2_SP_L3D3PHI3X2_L4D3PHI3X2_wr_en;
wire [5:0] SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3X2_L4D3PHI3X2(
.data_in(TE_L3D3PHI3X2_L4D3PHI3X2_SP_L3D3PHI3X2_L4D3PHI3X2),
.enable(TE_L3D3PHI3X2_L4D3PHI3X2_SP_L3D3PHI3X2_L4D3PHI3X2_wr_en),
.number_out(SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3),
.start(TE_L3D3PHI3X2_L4D3PHI3X2_start),
.done(SP_L3D3PHI3X2_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI3X2_L4D3PHI4X2_SP_L3D3PHI3X2_L4D3PHI4X2;
wire TE_L3D3PHI3X2_L4D3PHI4X2_SP_L3D3PHI3X2_L4D3PHI4X2_wr_en;
wire [5:0] SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3_number;
wire [8:0] SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3_read_add;
wire [11:0] SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3;
StubPairs  SP_L3D3PHI3X2_L4D3PHI4X2(
.data_in(TE_L3D3PHI3X2_L4D3PHI4X2_SP_L3D3PHI3X2_L4D3PHI4X2),
.enable(TE_L3D3PHI3X2_L4D3PHI4X2_SP_L3D3PHI3X2_L4D3PHI4X2_wr_en),
.number_out(SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3_number),
.read_add(SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3_read_add),
.data_out(SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3),
.start(TE_L3D3PHI3X2_L4D3PHI4X2_start),
.done(SP_L3D3PHI3X2_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L3D3_AS_L3D3n1;
wire VMR_L3D3_AS_L3D3n1_wr_en;
wire [10:0] AS_L3D3n1_TC_L3D3L4D3_read_add;
wire [35:0] AS_L3D3n1_TC_L3D3L4D3;
AllStubs  AS_L3D3n1(
.data_in(VMR_L3D3_AS_L3D3n1),
.enable(VMR_L3D3_AS_L3D3n1_wr_en),
.read_add(AS_L3D3n1_TC_L3D3L4D3_read_add),
.data_out(AS_L3D3n1_TC_L3D3L4D3),
.start(VMR_L3D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L4D3_AS_L4D3n1;
wire VMR_L4D3_AS_L4D3n1_wr_en;
wire [10:0] AS_L4D3n1_TC_L3D3L4D3_read_add;
wire [35:0] AS_L4D3n1_TC_L3D3L4D3;
AllStubs  AS_L4D3n1(
.data_in(VMR_L4D3_AS_L4D3n1),
.enable(VMR_L4D3_AS_L4D3n1_wr_en),
.read_add(AS_L4D3n1_TC_L3D3L4D3_read_add),
.data_out(AS_L4D3n1_TC_L3D3L4D3),
.start(VMR_L4D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI1X2_L4D4PHI1X1_SP_L3D3PHI1X2_L4D4PHI1X1;
wire TE_L3D3PHI1X2_L4D4PHI1X1_SP_L3D3PHI1X2_L4D4PHI1X1_wr_en;
wire [5:0] SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI1X2_L4D4PHI1X1(
.data_in(TE_L3D3PHI1X2_L4D4PHI1X1_SP_L3D3PHI1X2_L4D4PHI1X1),
.enable(TE_L3D3PHI1X2_L4D4PHI1X1_SP_L3D3PHI1X2_L4D4PHI1X1_wr_en),
.number_out(SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4),
.start(TE_L3D3PHI1X2_L4D4PHI1X1_start),
.done(SP_L3D3PHI1X2_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI1X2_L4D4PHI2X1_SP_L3D3PHI1X2_L4D4PHI2X1;
wire TE_L3D3PHI1X2_L4D4PHI2X1_SP_L3D3PHI1X2_L4D4PHI2X1_wr_en;
wire [5:0] SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI1X2_L4D4PHI2X1(
.data_in(TE_L3D3PHI1X2_L4D4PHI2X1_SP_L3D3PHI1X2_L4D4PHI2X1),
.enable(TE_L3D3PHI1X2_L4D4PHI2X1_SP_L3D3PHI1X2_L4D4PHI2X1_wr_en),
.number_out(SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4),
.start(TE_L3D3PHI1X2_L4D4PHI2X1_start),
.done(SP_L3D3PHI1X2_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI2X2_L4D4PHI2X1_SP_L3D3PHI2X2_L4D4PHI2X1;
wire TE_L3D3PHI2X2_L4D4PHI2X1_SP_L3D3PHI2X2_L4D4PHI2X1_wr_en;
wire [5:0] SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI2X2_L4D4PHI2X1(
.data_in(TE_L3D3PHI2X2_L4D4PHI2X1_SP_L3D3PHI2X2_L4D4PHI2X1),
.enable(TE_L3D3PHI2X2_L4D4PHI2X1_SP_L3D3PHI2X2_L4D4PHI2X1_wr_en),
.number_out(SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4),
.start(TE_L3D3PHI2X2_L4D4PHI2X1_start),
.done(SP_L3D3PHI2X2_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI2X2_L4D4PHI3X1_SP_L3D3PHI2X2_L4D4PHI3X1;
wire TE_L3D3PHI2X2_L4D4PHI3X1_SP_L3D3PHI2X2_L4D4PHI3X1_wr_en;
wire [5:0] SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI2X2_L4D4PHI3X1(
.data_in(TE_L3D3PHI2X2_L4D4PHI3X1_SP_L3D3PHI2X2_L4D4PHI3X1),
.enable(TE_L3D3PHI2X2_L4D4PHI3X1_SP_L3D3PHI2X2_L4D4PHI3X1_wr_en),
.number_out(SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4),
.start(TE_L3D3PHI2X2_L4D4PHI3X1_start),
.done(SP_L3D3PHI2X2_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI3X2_L4D4PHI3X1_SP_L3D3PHI3X2_L4D4PHI3X1;
wire TE_L3D3PHI3X2_L4D4PHI3X1_SP_L3D3PHI3X2_L4D4PHI3X1_wr_en;
wire [5:0] SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI3X2_L4D4PHI3X1(
.data_in(TE_L3D3PHI3X2_L4D4PHI3X1_SP_L3D3PHI3X2_L4D4PHI3X1),
.enable(TE_L3D3PHI3X2_L4D4PHI3X1_SP_L3D3PHI3X2_L4D4PHI3X1_wr_en),
.number_out(SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4),
.start(TE_L3D3PHI3X2_L4D4PHI3X1_start),
.done(SP_L3D3PHI3X2_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D3PHI3X2_L4D4PHI4X1_SP_L3D3PHI3X2_L4D4PHI4X1;
wire TE_L3D3PHI3X2_L4D4PHI4X1_SP_L3D3PHI3X2_L4D4PHI4X1_wr_en;
wire [5:0] SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4_number;
wire [8:0] SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4_read_add;
wire [11:0] SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4;
StubPairs  SP_L3D3PHI3X2_L4D4PHI4X1(
.data_in(TE_L3D3PHI3X2_L4D4PHI4X1_SP_L3D3PHI3X2_L4D4PHI4X1),
.enable(TE_L3D3PHI3X2_L4D4PHI4X1_SP_L3D3PHI3X2_L4D4PHI4X1_wr_en),
.number_out(SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4_number),
.read_add(SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4_read_add),
.data_out(SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4),
.start(TE_L3D3PHI3X2_L4D4PHI4X1_start),
.done(SP_L3D3PHI3X2_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L3D3_AS_L3D3n2;
wire VMR_L3D3_AS_L3D3n2_wr_en;
wire [10:0] AS_L3D3n2_TC_L3D3L4D4_read_add;
wire [35:0] AS_L3D3n2_TC_L3D3L4D4;
AllStubs  AS_L3D3n2(
.data_in(VMR_L3D3_AS_L3D3n2),
.enable(VMR_L3D3_AS_L3D3n2_wr_en),
.read_add(AS_L3D3n2_TC_L3D3L4D4_read_add),
.data_out(AS_L3D3n2_TC_L3D3L4D4),
.start(VMR_L3D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L4D4_AS_L4D4n1;
wire VMR_L4D4_AS_L4D4n1_wr_en;
wire [10:0] AS_L4D4n1_TC_L3D3L4D4_read_add;
wire [35:0] AS_L4D4n1_TC_L3D3L4D4;
AllStubs  AS_L4D4n1(
.data_in(VMR_L4D4_AS_L4D4n1),
.enable(VMR_L4D4_AS_L4D4n1_wr_en),
.read_add(AS_L4D4n1_TC_L3D3L4D4_read_add),
.data_out(AS_L4D4n1_TC_L3D3L4D4),
.start(VMR_L4D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI1X1_L4D4PHI1X1_SP_L3D4PHI1X1_L4D4PHI1X1;
wire TE_L3D4PHI1X1_L4D4PHI1X1_SP_L3D4PHI1X1_L4D4PHI1X1_wr_en;
wire [5:0] SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1X1_L4D4PHI1X1(
.data_in(TE_L3D4PHI1X1_L4D4PHI1X1_SP_L3D4PHI1X1_L4D4PHI1X1),
.enable(TE_L3D4PHI1X1_L4D4PHI1X1_SP_L3D4PHI1X1_L4D4PHI1X1_wr_en),
.number_out(SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4),
.start(TE_L3D4PHI1X1_L4D4PHI1X1_start),
.done(SP_L3D4PHI1X1_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI1X1_L4D4PHI2X1_SP_L3D4PHI1X1_L4D4PHI2X1;
wire TE_L3D4PHI1X1_L4D4PHI2X1_SP_L3D4PHI1X1_L4D4PHI2X1_wr_en;
wire [5:0] SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1X1_L4D4PHI2X1(
.data_in(TE_L3D4PHI1X1_L4D4PHI2X1_SP_L3D4PHI1X1_L4D4PHI2X1),
.enable(TE_L3D4PHI1X1_L4D4PHI2X1_SP_L3D4PHI1X1_L4D4PHI2X1_wr_en),
.number_out(SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4),
.start(TE_L3D4PHI1X1_L4D4PHI2X1_start),
.done(SP_L3D4PHI1X1_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI2X1_L4D4PHI2X1_SP_L3D4PHI2X1_L4D4PHI2X1;
wire TE_L3D4PHI2X1_L4D4PHI2X1_SP_L3D4PHI2X1_L4D4PHI2X1_wr_en;
wire [5:0] SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2X1_L4D4PHI2X1(
.data_in(TE_L3D4PHI2X1_L4D4PHI2X1_SP_L3D4PHI2X1_L4D4PHI2X1),
.enable(TE_L3D4PHI2X1_L4D4PHI2X1_SP_L3D4PHI2X1_L4D4PHI2X1_wr_en),
.number_out(SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4),
.start(TE_L3D4PHI2X1_L4D4PHI2X1_start),
.done(SP_L3D4PHI2X1_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI2X1_L4D4PHI3X1_SP_L3D4PHI2X1_L4D4PHI3X1;
wire TE_L3D4PHI2X1_L4D4PHI3X1_SP_L3D4PHI2X1_L4D4PHI3X1_wr_en;
wire [5:0] SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2X1_L4D4PHI3X1(
.data_in(TE_L3D4PHI2X1_L4D4PHI3X1_SP_L3D4PHI2X1_L4D4PHI3X1),
.enable(TE_L3D4PHI2X1_L4D4PHI3X1_SP_L3D4PHI2X1_L4D4PHI3X1_wr_en),
.number_out(SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4),
.start(TE_L3D4PHI2X1_L4D4PHI3X1_start),
.done(SP_L3D4PHI2X1_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI3X1_L4D4PHI3X1_SP_L3D4PHI3X1_L4D4PHI3X1;
wire TE_L3D4PHI3X1_L4D4PHI3X1_SP_L3D4PHI3X1_L4D4PHI3X1_wr_en;
wire [5:0] SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3X1_L4D4PHI3X1(
.data_in(TE_L3D4PHI3X1_L4D4PHI3X1_SP_L3D4PHI3X1_L4D4PHI3X1),
.enable(TE_L3D4PHI3X1_L4D4PHI3X1_SP_L3D4PHI3X1_L4D4PHI3X1_wr_en),
.number_out(SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4),
.start(TE_L3D4PHI3X1_L4D4PHI3X1_start),
.done(SP_L3D4PHI3X1_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI3X1_L4D4PHI4X1_SP_L3D4PHI3X1_L4D4PHI4X1;
wire TE_L3D4PHI3X1_L4D4PHI4X1_SP_L3D4PHI3X1_L4D4PHI4X1_wr_en;
wire [5:0] SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3X1_L4D4PHI4X1(
.data_in(TE_L3D4PHI3X1_L4D4PHI4X1_SP_L3D4PHI3X1_L4D4PHI4X1),
.enable(TE_L3D4PHI3X1_L4D4PHI4X1_SP_L3D4PHI3X1_L4D4PHI4X1_wr_en),
.number_out(SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4),
.start(TE_L3D4PHI3X1_L4D4PHI4X1_start),
.done(SP_L3D4PHI3X1_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI1X1_L4D4PHI1X2_SP_L3D4PHI1X1_L4D4PHI1X2;
wire TE_L3D4PHI1X1_L4D4PHI1X2_SP_L3D4PHI1X1_L4D4PHI1X2_wr_en;
wire [5:0] SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1X1_L4D4PHI1X2(
.data_in(TE_L3D4PHI1X1_L4D4PHI1X2_SP_L3D4PHI1X1_L4D4PHI1X2),
.enable(TE_L3D4PHI1X1_L4D4PHI1X2_SP_L3D4PHI1X1_L4D4PHI1X2_wr_en),
.number_out(SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4),
.start(TE_L3D4PHI1X1_L4D4PHI1X2_start),
.done(SP_L3D4PHI1X1_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI1X1_L4D4PHI2X2_SP_L3D4PHI1X1_L4D4PHI2X2;
wire TE_L3D4PHI1X1_L4D4PHI2X2_SP_L3D4PHI1X1_L4D4PHI2X2_wr_en;
wire [5:0] SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1X1_L4D4PHI2X2(
.data_in(TE_L3D4PHI1X1_L4D4PHI2X2_SP_L3D4PHI1X1_L4D4PHI2X2),
.enable(TE_L3D4PHI1X1_L4D4PHI2X2_SP_L3D4PHI1X1_L4D4PHI2X2_wr_en),
.number_out(SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4),
.start(TE_L3D4PHI1X1_L4D4PHI2X2_start),
.done(SP_L3D4PHI1X1_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI2X1_L4D4PHI2X2_SP_L3D4PHI2X1_L4D4PHI2X2;
wire TE_L3D4PHI2X1_L4D4PHI2X2_SP_L3D4PHI2X1_L4D4PHI2X2_wr_en;
wire [5:0] SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2X1_L4D4PHI2X2(
.data_in(TE_L3D4PHI2X1_L4D4PHI2X2_SP_L3D4PHI2X1_L4D4PHI2X2),
.enable(TE_L3D4PHI2X1_L4D4PHI2X2_SP_L3D4PHI2X1_L4D4PHI2X2_wr_en),
.number_out(SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4),
.start(TE_L3D4PHI2X1_L4D4PHI2X2_start),
.done(SP_L3D4PHI2X1_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI2X1_L4D4PHI3X2_SP_L3D4PHI2X1_L4D4PHI3X2;
wire TE_L3D4PHI2X1_L4D4PHI3X2_SP_L3D4PHI2X1_L4D4PHI3X2_wr_en;
wire [5:0] SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2X1_L4D4PHI3X2(
.data_in(TE_L3D4PHI2X1_L4D4PHI3X2_SP_L3D4PHI2X1_L4D4PHI3X2),
.enable(TE_L3D4PHI2X1_L4D4PHI3X2_SP_L3D4PHI2X1_L4D4PHI3X2_wr_en),
.number_out(SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4),
.start(TE_L3D4PHI2X1_L4D4PHI3X2_start),
.done(SP_L3D4PHI2X1_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI3X1_L4D4PHI3X2_SP_L3D4PHI3X1_L4D4PHI3X2;
wire TE_L3D4PHI3X1_L4D4PHI3X2_SP_L3D4PHI3X1_L4D4PHI3X2_wr_en;
wire [5:0] SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3X1_L4D4PHI3X2(
.data_in(TE_L3D4PHI3X1_L4D4PHI3X2_SP_L3D4PHI3X1_L4D4PHI3X2),
.enable(TE_L3D4PHI3X1_L4D4PHI3X2_SP_L3D4PHI3X1_L4D4PHI3X2_wr_en),
.number_out(SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4),
.start(TE_L3D4PHI3X1_L4D4PHI3X2_start),
.done(SP_L3D4PHI3X1_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI3X1_L4D4PHI4X2_SP_L3D4PHI3X1_L4D4PHI4X2;
wire TE_L3D4PHI3X1_L4D4PHI4X2_SP_L3D4PHI3X1_L4D4PHI4X2_wr_en;
wire [5:0] SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3X1_L4D4PHI4X2(
.data_in(TE_L3D4PHI3X1_L4D4PHI4X2_SP_L3D4PHI3X1_L4D4PHI4X2),
.enable(TE_L3D4PHI3X1_L4D4PHI4X2_SP_L3D4PHI3X1_L4D4PHI4X2_wr_en),
.number_out(SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4),
.start(TE_L3D4PHI3X1_L4D4PHI4X2_start),
.done(SP_L3D4PHI3X1_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI1X2_L4D4PHI1X2_SP_L3D4PHI1X2_L4D4PHI1X2;
wire TE_L3D4PHI1X2_L4D4PHI1X2_SP_L3D4PHI1X2_L4D4PHI1X2_wr_en;
wire [5:0] SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1X2_L4D4PHI1X2(
.data_in(TE_L3D4PHI1X2_L4D4PHI1X2_SP_L3D4PHI1X2_L4D4PHI1X2),
.enable(TE_L3D4PHI1X2_L4D4PHI1X2_SP_L3D4PHI1X2_L4D4PHI1X2_wr_en),
.number_out(SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4),
.start(TE_L3D4PHI1X2_L4D4PHI1X2_start),
.done(SP_L3D4PHI1X2_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI1X2_L4D4PHI2X2_SP_L3D4PHI1X2_L4D4PHI2X2;
wire TE_L3D4PHI1X2_L4D4PHI2X2_SP_L3D4PHI1X2_L4D4PHI2X2_wr_en;
wire [5:0] SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI1X2_L4D4PHI2X2(
.data_in(TE_L3D4PHI1X2_L4D4PHI2X2_SP_L3D4PHI1X2_L4D4PHI2X2),
.enable(TE_L3D4PHI1X2_L4D4PHI2X2_SP_L3D4PHI1X2_L4D4PHI2X2_wr_en),
.number_out(SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4),
.start(TE_L3D4PHI1X2_L4D4PHI2X2_start),
.done(SP_L3D4PHI1X2_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI2X2_L4D4PHI2X2_SP_L3D4PHI2X2_L4D4PHI2X2;
wire TE_L3D4PHI2X2_L4D4PHI2X2_SP_L3D4PHI2X2_L4D4PHI2X2_wr_en;
wire [5:0] SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2X2_L4D4PHI2X2(
.data_in(TE_L3D4PHI2X2_L4D4PHI2X2_SP_L3D4PHI2X2_L4D4PHI2X2),
.enable(TE_L3D4PHI2X2_L4D4PHI2X2_SP_L3D4PHI2X2_L4D4PHI2X2_wr_en),
.number_out(SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4),
.start(TE_L3D4PHI2X2_L4D4PHI2X2_start),
.done(SP_L3D4PHI2X2_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI2X2_L4D4PHI3X2_SP_L3D4PHI2X2_L4D4PHI3X2;
wire TE_L3D4PHI2X2_L4D4PHI3X2_SP_L3D4PHI2X2_L4D4PHI3X2_wr_en;
wire [5:0] SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI2X2_L4D4PHI3X2(
.data_in(TE_L3D4PHI2X2_L4D4PHI3X2_SP_L3D4PHI2X2_L4D4PHI3X2),
.enable(TE_L3D4PHI2X2_L4D4PHI3X2_SP_L3D4PHI2X2_L4D4PHI3X2_wr_en),
.number_out(SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4),
.start(TE_L3D4PHI2X2_L4D4PHI3X2_start),
.done(SP_L3D4PHI2X2_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI3X2_L4D4PHI3X2_SP_L3D4PHI3X2_L4D4PHI3X2;
wire TE_L3D4PHI3X2_L4D4PHI3X2_SP_L3D4PHI3X2_L4D4PHI3X2_wr_en;
wire [5:0] SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3X2_L4D4PHI3X2(
.data_in(TE_L3D4PHI3X2_L4D4PHI3X2_SP_L3D4PHI3X2_L4D4PHI3X2),
.enable(TE_L3D4PHI3X2_L4D4PHI3X2_SP_L3D4PHI3X2_L4D4PHI3X2_wr_en),
.number_out(SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4),
.start(TE_L3D4PHI3X2_L4D4PHI3X2_start),
.done(SP_L3D4PHI3X2_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L3D4PHI3X2_L4D4PHI4X2_SP_L3D4PHI3X2_L4D4PHI4X2;
wire TE_L3D4PHI3X2_L4D4PHI4X2_SP_L3D4PHI3X2_L4D4PHI4X2_wr_en;
wire [5:0] SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4_number;
wire [8:0] SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4_read_add;
wire [11:0] SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4;
StubPairs  SP_L3D4PHI3X2_L4D4PHI4X2(
.data_in(TE_L3D4PHI3X2_L4D4PHI4X2_SP_L3D4PHI3X2_L4D4PHI4X2),
.enable(TE_L3D4PHI3X2_L4D4PHI4X2_SP_L3D4PHI3X2_L4D4PHI4X2_wr_en),
.number_out(SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4_number),
.read_add(SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4_read_add),
.data_out(SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4),
.start(TE_L3D4PHI3X2_L4D4PHI4X2_start),
.done(SP_L3D4PHI3X2_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L3D4_AS_L3D4n1;
wire VMR_L3D4_AS_L3D4n1_wr_en;
wire [10:0] AS_L3D4n1_TC_L3D4L4D4_read_add;
wire [35:0] AS_L3D4n1_TC_L3D4L4D4;
AllStubs  AS_L3D4n1(
.data_in(VMR_L3D4_AS_L3D4n1),
.enable(VMR_L3D4_AS_L3D4n1_wr_en),
.read_add(AS_L3D4n1_TC_L3D4L4D4_read_add),
.data_out(AS_L3D4n1_TC_L3D4L4D4),
.start(VMR_L3D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L4D4_AS_L4D4n2;
wire VMR_L4D4_AS_L4D4n2_wr_en;
wire [10:0] AS_L4D4n2_TC_L3D4L4D4_read_add;
wire [35:0] AS_L4D4n2_TC_L3D4L4D4;
AllStubs  AS_L4D4n2(
.data_in(VMR_L4D4_AS_L4D4n2),
.enable(VMR_L4D4_AS_L4D4n2_wr_en),
.read_add(AS_L4D4n2_TC_L3D4L4D4_read_add),
.data_out(AS_L4D4n2_TC_L3D4L4D4),
.start(VMR_L4D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI1X1_L6D3PHI1X1_SP_L5D3PHI1X1_L6D3PHI1X1;
wire TE_L5D3PHI1X1_L6D3PHI1X1_SP_L5D3PHI1X1_L6D3PHI1X1_wr_en;
wire [5:0] SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1X1_L6D3PHI1X1(
.data_in(TE_L5D3PHI1X1_L6D3PHI1X1_SP_L5D3PHI1X1_L6D3PHI1X1),
.enable(TE_L5D3PHI1X1_L6D3PHI1X1_SP_L5D3PHI1X1_L6D3PHI1X1_wr_en),
.number_out(SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3),
.start(TE_L5D3PHI1X1_L6D3PHI1X1_start),
.done(SP_L5D3PHI1X1_L6D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI1X1_L6D3PHI2X1_SP_L5D3PHI1X1_L6D3PHI2X1;
wire TE_L5D3PHI1X1_L6D3PHI2X1_SP_L5D3PHI1X1_L6D3PHI2X1_wr_en;
wire [5:0] SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1X1_L6D3PHI2X1(
.data_in(TE_L5D3PHI1X1_L6D3PHI2X1_SP_L5D3PHI1X1_L6D3PHI2X1),
.enable(TE_L5D3PHI1X1_L6D3PHI2X1_SP_L5D3PHI1X1_L6D3PHI2X1_wr_en),
.number_out(SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3),
.start(TE_L5D3PHI1X1_L6D3PHI2X1_start),
.done(SP_L5D3PHI1X1_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI2X1_L6D3PHI2X1_SP_L5D3PHI2X1_L6D3PHI2X1;
wire TE_L5D3PHI2X1_L6D3PHI2X1_SP_L5D3PHI2X1_L6D3PHI2X1_wr_en;
wire [5:0] SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2X1_L6D3PHI2X1(
.data_in(TE_L5D3PHI2X1_L6D3PHI2X1_SP_L5D3PHI2X1_L6D3PHI2X1),
.enable(TE_L5D3PHI2X1_L6D3PHI2X1_SP_L5D3PHI2X1_L6D3PHI2X1_wr_en),
.number_out(SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3),
.start(TE_L5D3PHI2X1_L6D3PHI2X1_start),
.done(SP_L5D3PHI2X1_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI2X1_L6D3PHI3X1_SP_L5D3PHI2X1_L6D3PHI3X1;
wire TE_L5D3PHI2X1_L6D3PHI3X1_SP_L5D3PHI2X1_L6D3PHI3X1_wr_en;
wire [5:0] SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2X1_L6D3PHI3X1(
.data_in(TE_L5D3PHI2X1_L6D3PHI3X1_SP_L5D3PHI2X1_L6D3PHI3X1),
.enable(TE_L5D3PHI2X1_L6D3PHI3X1_SP_L5D3PHI2X1_L6D3PHI3X1_wr_en),
.number_out(SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3),
.start(TE_L5D3PHI2X1_L6D3PHI3X1_start),
.done(SP_L5D3PHI2X1_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI3X1_L6D3PHI3X1_SP_L5D3PHI3X1_L6D3PHI3X1;
wire TE_L5D3PHI3X1_L6D3PHI3X1_SP_L5D3PHI3X1_L6D3PHI3X1_wr_en;
wire [5:0] SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3X1_L6D3PHI3X1(
.data_in(TE_L5D3PHI3X1_L6D3PHI3X1_SP_L5D3PHI3X1_L6D3PHI3X1),
.enable(TE_L5D3PHI3X1_L6D3PHI3X1_SP_L5D3PHI3X1_L6D3PHI3X1_wr_en),
.number_out(SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3),
.start(TE_L5D3PHI3X1_L6D3PHI3X1_start),
.done(SP_L5D3PHI3X1_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI3X1_L6D3PHI4X1_SP_L5D3PHI3X1_L6D3PHI4X1;
wire TE_L5D3PHI3X1_L6D3PHI4X1_SP_L5D3PHI3X1_L6D3PHI4X1_wr_en;
wire [5:0] SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3X1_L6D3PHI4X1(
.data_in(TE_L5D3PHI3X1_L6D3PHI4X1_SP_L5D3PHI3X1_L6D3PHI4X1),
.enable(TE_L5D3PHI3X1_L6D3PHI4X1_SP_L5D3PHI3X1_L6D3PHI4X1_wr_en),
.number_out(SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3),
.start(TE_L5D3PHI3X1_L6D3PHI4X1_start),
.done(SP_L5D3PHI3X1_L6D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI1X1_L6D3PHI1X2_SP_L5D3PHI1X1_L6D3PHI1X2;
wire TE_L5D3PHI1X1_L6D3PHI1X2_SP_L5D3PHI1X1_L6D3PHI1X2_wr_en;
wire [5:0] SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1X1_L6D3PHI1X2(
.data_in(TE_L5D3PHI1X1_L6D3PHI1X2_SP_L5D3PHI1X1_L6D3PHI1X2),
.enable(TE_L5D3PHI1X1_L6D3PHI1X2_SP_L5D3PHI1X1_L6D3PHI1X2_wr_en),
.number_out(SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3),
.start(TE_L5D3PHI1X1_L6D3PHI1X2_start),
.done(SP_L5D3PHI1X1_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI1X1_L6D3PHI2X2_SP_L5D3PHI1X1_L6D3PHI2X2;
wire TE_L5D3PHI1X1_L6D3PHI2X2_SP_L5D3PHI1X1_L6D3PHI2X2_wr_en;
wire [5:0] SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1X1_L6D3PHI2X2(
.data_in(TE_L5D3PHI1X1_L6D3PHI2X2_SP_L5D3PHI1X1_L6D3PHI2X2),
.enable(TE_L5D3PHI1X1_L6D3PHI2X2_SP_L5D3PHI1X1_L6D3PHI2X2_wr_en),
.number_out(SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3),
.start(TE_L5D3PHI1X1_L6D3PHI2X2_start),
.done(SP_L5D3PHI1X1_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI2X1_L6D3PHI2X2_SP_L5D3PHI2X1_L6D3PHI2X2;
wire TE_L5D3PHI2X1_L6D3PHI2X2_SP_L5D3PHI2X1_L6D3PHI2X2_wr_en;
wire [5:0] SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2X1_L6D3PHI2X2(
.data_in(TE_L5D3PHI2X1_L6D3PHI2X2_SP_L5D3PHI2X1_L6D3PHI2X2),
.enable(TE_L5D3PHI2X1_L6D3PHI2X2_SP_L5D3PHI2X1_L6D3PHI2X2_wr_en),
.number_out(SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3),
.start(TE_L5D3PHI2X1_L6D3PHI2X2_start),
.done(SP_L5D3PHI2X1_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI2X1_L6D3PHI3X2_SP_L5D3PHI2X1_L6D3PHI3X2;
wire TE_L5D3PHI2X1_L6D3PHI3X2_SP_L5D3PHI2X1_L6D3PHI3X2_wr_en;
wire [5:0] SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2X1_L6D3PHI3X2(
.data_in(TE_L5D3PHI2X1_L6D3PHI3X2_SP_L5D3PHI2X1_L6D3PHI3X2),
.enable(TE_L5D3PHI2X1_L6D3PHI3X2_SP_L5D3PHI2X1_L6D3PHI3X2_wr_en),
.number_out(SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3),
.start(TE_L5D3PHI2X1_L6D3PHI3X2_start),
.done(SP_L5D3PHI2X1_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI3X1_L6D3PHI3X2_SP_L5D3PHI3X1_L6D3PHI3X2;
wire TE_L5D3PHI3X1_L6D3PHI3X2_SP_L5D3PHI3X1_L6D3PHI3X2_wr_en;
wire [5:0] SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3X1_L6D3PHI3X2(
.data_in(TE_L5D3PHI3X1_L6D3PHI3X2_SP_L5D3PHI3X1_L6D3PHI3X2),
.enable(TE_L5D3PHI3X1_L6D3PHI3X2_SP_L5D3PHI3X1_L6D3PHI3X2_wr_en),
.number_out(SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3),
.start(TE_L5D3PHI3X1_L6D3PHI3X2_start),
.done(SP_L5D3PHI3X1_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI3X1_L6D3PHI4X2_SP_L5D3PHI3X1_L6D3PHI4X2;
wire TE_L5D3PHI3X1_L6D3PHI4X2_SP_L5D3PHI3X1_L6D3PHI4X2_wr_en;
wire [5:0] SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3X1_L6D3PHI4X2(
.data_in(TE_L5D3PHI3X1_L6D3PHI4X2_SP_L5D3PHI3X1_L6D3PHI4X2),
.enable(TE_L5D3PHI3X1_L6D3PHI4X2_SP_L5D3PHI3X1_L6D3PHI4X2_wr_en),
.number_out(SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3),
.start(TE_L5D3PHI3X1_L6D3PHI4X2_start),
.done(SP_L5D3PHI3X1_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI1X2_L6D3PHI1X2_SP_L5D3PHI1X2_L6D3PHI1X2;
wire TE_L5D3PHI1X2_L6D3PHI1X2_SP_L5D3PHI1X2_L6D3PHI1X2_wr_en;
wire [5:0] SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1X2_L6D3PHI1X2(
.data_in(TE_L5D3PHI1X2_L6D3PHI1X2_SP_L5D3PHI1X2_L6D3PHI1X2),
.enable(TE_L5D3PHI1X2_L6D3PHI1X2_SP_L5D3PHI1X2_L6D3PHI1X2_wr_en),
.number_out(SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3),
.start(TE_L5D3PHI1X2_L6D3PHI1X2_start),
.done(SP_L5D3PHI1X2_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI1X2_L6D3PHI2X2_SP_L5D3PHI1X2_L6D3PHI2X2;
wire TE_L5D3PHI1X2_L6D3PHI2X2_SP_L5D3PHI1X2_L6D3PHI2X2_wr_en;
wire [5:0] SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI1X2_L6D3PHI2X2(
.data_in(TE_L5D3PHI1X2_L6D3PHI2X2_SP_L5D3PHI1X2_L6D3PHI2X2),
.enable(TE_L5D3PHI1X2_L6D3PHI2X2_SP_L5D3PHI1X2_L6D3PHI2X2_wr_en),
.number_out(SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3),
.start(TE_L5D3PHI1X2_L6D3PHI2X2_start),
.done(SP_L5D3PHI1X2_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI2X2_L6D3PHI2X2_SP_L5D3PHI2X2_L6D3PHI2X2;
wire TE_L5D3PHI2X2_L6D3PHI2X2_SP_L5D3PHI2X2_L6D3PHI2X2_wr_en;
wire [5:0] SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2X2_L6D3PHI2X2(
.data_in(TE_L5D3PHI2X2_L6D3PHI2X2_SP_L5D3PHI2X2_L6D3PHI2X2),
.enable(TE_L5D3PHI2X2_L6D3PHI2X2_SP_L5D3PHI2X2_L6D3PHI2X2_wr_en),
.number_out(SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3),
.start(TE_L5D3PHI2X2_L6D3PHI2X2_start),
.done(SP_L5D3PHI2X2_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI2X2_L6D3PHI3X2_SP_L5D3PHI2X2_L6D3PHI3X2;
wire TE_L5D3PHI2X2_L6D3PHI3X2_SP_L5D3PHI2X2_L6D3PHI3X2_wr_en;
wire [5:0] SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI2X2_L6D3PHI3X2(
.data_in(TE_L5D3PHI2X2_L6D3PHI3X2_SP_L5D3PHI2X2_L6D3PHI3X2),
.enable(TE_L5D3PHI2X2_L6D3PHI3X2_SP_L5D3PHI2X2_L6D3PHI3X2_wr_en),
.number_out(SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3),
.start(TE_L5D3PHI2X2_L6D3PHI3X2_start),
.done(SP_L5D3PHI2X2_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI3X2_L6D3PHI3X2_SP_L5D3PHI3X2_L6D3PHI3X2;
wire TE_L5D3PHI3X2_L6D3PHI3X2_SP_L5D3PHI3X2_L6D3PHI3X2_wr_en;
wire [5:0] SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3X2_L6D3PHI3X2(
.data_in(TE_L5D3PHI3X2_L6D3PHI3X2_SP_L5D3PHI3X2_L6D3PHI3X2),
.enable(TE_L5D3PHI3X2_L6D3PHI3X2_SP_L5D3PHI3X2_L6D3PHI3X2_wr_en),
.number_out(SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3),
.start(TE_L5D3PHI3X2_L6D3PHI3X2_start),
.done(SP_L5D3PHI3X2_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI3X2_L6D3PHI4X2_SP_L5D3PHI3X2_L6D3PHI4X2;
wire TE_L5D3PHI3X2_L6D3PHI4X2_SP_L5D3PHI3X2_L6D3PHI4X2_wr_en;
wire [5:0] SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3_number;
wire [8:0] SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3_read_add;
wire [11:0] SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3;
StubPairs  SP_L5D3PHI3X2_L6D3PHI4X2(
.data_in(TE_L5D3PHI3X2_L6D3PHI4X2_SP_L5D3PHI3X2_L6D3PHI4X2),
.enable(TE_L5D3PHI3X2_L6D3PHI4X2_SP_L5D3PHI3X2_L6D3PHI4X2_wr_en),
.number_out(SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3_number),
.read_add(SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3_read_add),
.data_out(SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3),
.start(TE_L5D3PHI3X2_L6D3PHI4X2_start),
.done(SP_L5D3PHI3X2_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L5D3_AS_L5D3n1;
wire VMR_L5D3_AS_L5D3n1_wr_en;
wire [10:0] AS_L5D3n1_TC_L5D3L6D3_read_add;
wire [35:0] AS_L5D3n1_TC_L5D3L6D3;
AllStubs  AS_L5D3n1(
.data_in(VMR_L5D3_AS_L5D3n1),
.enable(VMR_L5D3_AS_L5D3n1_wr_en),
.read_add(AS_L5D3n1_TC_L5D3L6D3_read_add),
.data_out(AS_L5D3n1_TC_L5D3L6D3),
.start(VMR_L5D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L6D3_AS_L6D3n1;
wire VMR_L6D3_AS_L6D3n1_wr_en;
wire [10:0] AS_L6D3n1_TC_L5D3L6D3_read_add;
wire [35:0] AS_L6D3n1_TC_L5D3L6D3;
AllStubs  AS_L6D3n1(
.data_in(VMR_L6D3_AS_L6D3n1),
.enable(VMR_L6D3_AS_L6D3n1_wr_en),
.read_add(AS_L6D3n1_TC_L5D3L6D3_read_add),
.data_out(AS_L6D3n1_TC_L5D3L6D3),
.start(VMR_L6D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI1X2_L6D4PHI1X1_SP_L5D3PHI1X2_L6D4PHI1X1;
wire TE_L5D3PHI1X2_L6D4PHI1X1_SP_L5D3PHI1X2_L6D4PHI1X1_wr_en;
wire [5:0] SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI1X2_L6D4PHI1X1(
.data_in(TE_L5D3PHI1X2_L6D4PHI1X1_SP_L5D3PHI1X2_L6D4PHI1X1),
.enable(TE_L5D3PHI1X2_L6D4PHI1X1_SP_L5D3PHI1X2_L6D4PHI1X1_wr_en),
.number_out(SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4),
.start(TE_L5D3PHI1X2_L6D4PHI1X1_start),
.done(SP_L5D3PHI1X2_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI1X2_L6D4PHI2X1_SP_L5D3PHI1X2_L6D4PHI2X1;
wire TE_L5D3PHI1X2_L6D4PHI2X1_SP_L5D3PHI1X2_L6D4PHI2X1_wr_en;
wire [5:0] SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI1X2_L6D4PHI2X1(
.data_in(TE_L5D3PHI1X2_L6D4PHI2X1_SP_L5D3PHI1X2_L6D4PHI2X1),
.enable(TE_L5D3PHI1X2_L6D4PHI2X1_SP_L5D3PHI1X2_L6D4PHI2X1_wr_en),
.number_out(SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4),
.start(TE_L5D3PHI1X2_L6D4PHI2X1_start),
.done(SP_L5D3PHI1X2_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI2X2_L6D4PHI2X1_SP_L5D3PHI2X2_L6D4PHI2X1;
wire TE_L5D3PHI2X2_L6D4PHI2X1_SP_L5D3PHI2X2_L6D4PHI2X1_wr_en;
wire [5:0] SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI2X2_L6D4PHI2X1(
.data_in(TE_L5D3PHI2X2_L6D4PHI2X1_SP_L5D3PHI2X2_L6D4PHI2X1),
.enable(TE_L5D3PHI2X2_L6D4PHI2X1_SP_L5D3PHI2X2_L6D4PHI2X1_wr_en),
.number_out(SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4),
.start(TE_L5D3PHI2X2_L6D4PHI2X1_start),
.done(SP_L5D3PHI2X2_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI2X2_L6D4PHI3X1_SP_L5D3PHI2X2_L6D4PHI3X1;
wire TE_L5D3PHI2X2_L6D4PHI3X1_SP_L5D3PHI2X2_L6D4PHI3X1_wr_en;
wire [5:0] SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI2X2_L6D4PHI3X1(
.data_in(TE_L5D3PHI2X2_L6D4PHI3X1_SP_L5D3PHI2X2_L6D4PHI3X1),
.enable(TE_L5D3PHI2X2_L6D4PHI3X1_SP_L5D3PHI2X2_L6D4PHI3X1_wr_en),
.number_out(SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4),
.start(TE_L5D3PHI2X2_L6D4PHI3X1_start),
.done(SP_L5D3PHI2X2_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI3X2_L6D4PHI3X1_SP_L5D3PHI3X2_L6D4PHI3X1;
wire TE_L5D3PHI3X2_L6D4PHI3X1_SP_L5D3PHI3X2_L6D4PHI3X1_wr_en;
wire [5:0] SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI3X2_L6D4PHI3X1(
.data_in(TE_L5D3PHI3X2_L6D4PHI3X1_SP_L5D3PHI3X2_L6D4PHI3X1),
.enable(TE_L5D3PHI3X2_L6D4PHI3X1_SP_L5D3PHI3X2_L6D4PHI3X1_wr_en),
.number_out(SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4),
.start(TE_L5D3PHI3X2_L6D4PHI3X1_start),
.done(SP_L5D3PHI3X2_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D3PHI3X2_L6D4PHI4X1_SP_L5D3PHI3X2_L6D4PHI4X1;
wire TE_L5D3PHI3X2_L6D4PHI4X1_SP_L5D3PHI3X2_L6D4PHI4X1_wr_en;
wire [5:0] SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4_number;
wire [8:0] SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4_read_add;
wire [11:0] SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4;
StubPairs  SP_L5D3PHI3X2_L6D4PHI4X1(
.data_in(TE_L5D3PHI3X2_L6D4PHI4X1_SP_L5D3PHI3X2_L6D4PHI4X1),
.enable(TE_L5D3PHI3X2_L6D4PHI4X1_SP_L5D3PHI3X2_L6D4PHI4X1_wr_en),
.number_out(SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4_number),
.read_add(SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4_read_add),
.data_out(SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4),
.start(TE_L5D3PHI3X2_L6D4PHI4X1_start),
.done(SP_L5D3PHI3X2_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L5D3_AS_L5D3n2;
wire VMR_L5D3_AS_L5D3n2_wr_en;
wire [10:0] AS_L5D3n2_TC_L5D3L6D4_read_add;
wire [35:0] AS_L5D3n2_TC_L5D3L6D4;
AllStubs  AS_L5D3n2(
.data_in(VMR_L5D3_AS_L5D3n2),
.enable(VMR_L5D3_AS_L5D3n2_wr_en),
.read_add(AS_L5D3n2_TC_L5D3L6D4_read_add),
.data_out(AS_L5D3n2_TC_L5D3L6D4),
.start(VMR_L5D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L6D4_AS_L6D4n1;
wire VMR_L6D4_AS_L6D4n1_wr_en;
wire [10:0] AS_L6D4n1_TC_L5D3L6D4_read_add;
wire [35:0] AS_L6D4n1_TC_L5D3L6D4;
AllStubs  AS_L6D4n1(
.data_in(VMR_L6D4_AS_L6D4n1),
.enable(VMR_L6D4_AS_L6D4n1_wr_en),
.read_add(AS_L6D4n1_TC_L5D3L6D4_read_add),
.data_out(AS_L6D4n1_TC_L5D3L6D4),
.start(VMR_L6D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI1X1_L6D4PHI1X1_SP_L5D4PHI1X1_L6D4PHI1X1;
wire TE_L5D4PHI1X1_L6D4PHI1X1_SP_L5D4PHI1X1_L6D4PHI1X1_wr_en;
wire [5:0] SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1X1_L6D4PHI1X1(
.data_in(TE_L5D4PHI1X1_L6D4PHI1X1_SP_L5D4PHI1X1_L6D4PHI1X1),
.enable(TE_L5D4PHI1X1_L6D4PHI1X1_SP_L5D4PHI1X1_L6D4PHI1X1_wr_en),
.number_out(SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4),
.start(TE_L5D4PHI1X1_L6D4PHI1X1_start),
.done(SP_L5D4PHI1X1_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI1X1_L6D4PHI2X1_SP_L5D4PHI1X1_L6D4PHI2X1;
wire TE_L5D4PHI1X1_L6D4PHI2X1_SP_L5D4PHI1X1_L6D4PHI2X1_wr_en;
wire [5:0] SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1X1_L6D4PHI2X1(
.data_in(TE_L5D4PHI1X1_L6D4PHI2X1_SP_L5D4PHI1X1_L6D4PHI2X1),
.enable(TE_L5D4PHI1X1_L6D4PHI2X1_SP_L5D4PHI1X1_L6D4PHI2X1_wr_en),
.number_out(SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4),
.start(TE_L5D4PHI1X1_L6D4PHI2X1_start),
.done(SP_L5D4PHI1X1_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI2X1_L6D4PHI2X1_SP_L5D4PHI2X1_L6D4PHI2X1;
wire TE_L5D4PHI2X1_L6D4PHI2X1_SP_L5D4PHI2X1_L6D4PHI2X1_wr_en;
wire [5:0] SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2X1_L6D4PHI2X1(
.data_in(TE_L5D4PHI2X1_L6D4PHI2X1_SP_L5D4PHI2X1_L6D4PHI2X1),
.enable(TE_L5D4PHI2X1_L6D4PHI2X1_SP_L5D4PHI2X1_L6D4PHI2X1_wr_en),
.number_out(SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4),
.start(TE_L5D4PHI2X1_L6D4PHI2X1_start),
.done(SP_L5D4PHI2X1_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI2X1_L6D4PHI3X1_SP_L5D4PHI2X1_L6D4PHI3X1;
wire TE_L5D4PHI2X1_L6D4PHI3X1_SP_L5D4PHI2X1_L6D4PHI3X1_wr_en;
wire [5:0] SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2X1_L6D4PHI3X1(
.data_in(TE_L5D4PHI2X1_L6D4PHI3X1_SP_L5D4PHI2X1_L6D4PHI3X1),
.enable(TE_L5D4PHI2X1_L6D4PHI3X1_SP_L5D4PHI2X1_L6D4PHI3X1_wr_en),
.number_out(SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4),
.start(TE_L5D4PHI2X1_L6D4PHI3X1_start),
.done(SP_L5D4PHI2X1_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI3X1_L6D4PHI3X1_SP_L5D4PHI3X1_L6D4PHI3X1;
wire TE_L5D4PHI3X1_L6D4PHI3X1_SP_L5D4PHI3X1_L6D4PHI3X1_wr_en;
wire [5:0] SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3X1_L6D4PHI3X1(
.data_in(TE_L5D4PHI3X1_L6D4PHI3X1_SP_L5D4PHI3X1_L6D4PHI3X1),
.enable(TE_L5D4PHI3X1_L6D4PHI3X1_SP_L5D4PHI3X1_L6D4PHI3X1_wr_en),
.number_out(SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4),
.start(TE_L5D4PHI3X1_L6D4PHI3X1_start),
.done(SP_L5D4PHI3X1_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI3X1_L6D4PHI4X1_SP_L5D4PHI3X1_L6D4PHI4X1;
wire TE_L5D4PHI3X1_L6D4PHI4X1_SP_L5D4PHI3X1_L6D4PHI4X1_wr_en;
wire [5:0] SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3X1_L6D4PHI4X1(
.data_in(TE_L5D4PHI3X1_L6D4PHI4X1_SP_L5D4PHI3X1_L6D4PHI4X1),
.enable(TE_L5D4PHI3X1_L6D4PHI4X1_SP_L5D4PHI3X1_L6D4PHI4X1_wr_en),
.number_out(SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4),
.start(TE_L5D4PHI3X1_L6D4PHI4X1_start),
.done(SP_L5D4PHI3X1_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI1X1_L6D4PHI1X2_SP_L5D4PHI1X1_L6D4PHI1X2;
wire TE_L5D4PHI1X1_L6D4PHI1X2_SP_L5D4PHI1X1_L6D4PHI1X2_wr_en;
wire [5:0] SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1X1_L6D4PHI1X2(
.data_in(TE_L5D4PHI1X1_L6D4PHI1X2_SP_L5D4PHI1X1_L6D4PHI1X2),
.enable(TE_L5D4PHI1X1_L6D4PHI1X2_SP_L5D4PHI1X1_L6D4PHI1X2_wr_en),
.number_out(SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4),
.start(TE_L5D4PHI1X1_L6D4PHI1X2_start),
.done(SP_L5D4PHI1X1_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI1X1_L6D4PHI2X2_SP_L5D4PHI1X1_L6D4PHI2X2;
wire TE_L5D4PHI1X1_L6D4PHI2X2_SP_L5D4PHI1X1_L6D4PHI2X2_wr_en;
wire [5:0] SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1X1_L6D4PHI2X2(
.data_in(TE_L5D4PHI1X1_L6D4PHI2X2_SP_L5D4PHI1X1_L6D4PHI2X2),
.enable(TE_L5D4PHI1X1_L6D4PHI2X2_SP_L5D4PHI1X1_L6D4PHI2X2_wr_en),
.number_out(SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4),
.start(TE_L5D4PHI1X1_L6D4PHI2X2_start),
.done(SP_L5D4PHI1X1_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI2X1_L6D4PHI2X2_SP_L5D4PHI2X1_L6D4PHI2X2;
wire TE_L5D4PHI2X1_L6D4PHI2X2_SP_L5D4PHI2X1_L6D4PHI2X2_wr_en;
wire [5:0] SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2X1_L6D4PHI2X2(
.data_in(TE_L5D4PHI2X1_L6D4PHI2X2_SP_L5D4PHI2X1_L6D4PHI2X2),
.enable(TE_L5D4PHI2X1_L6D4PHI2X2_SP_L5D4PHI2X1_L6D4PHI2X2_wr_en),
.number_out(SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4),
.start(TE_L5D4PHI2X1_L6D4PHI2X2_start),
.done(SP_L5D4PHI2X1_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI2X1_L6D4PHI3X2_SP_L5D4PHI2X1_L6D4PHI3X2;
wire TE_L5D4PHI2X1_L6D4PHI3X2_SP_L5D4PHI2X1_L6D4PHI3X2_wr_en;
wire [5:0] SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2X1_L6D4PHI3X2(
.data_in(TE_L5D4PHI2X1_L6D4PHI3X2_SP_L5D4PHI2X1_L6D4PHI3X2),
.enable(TE_L5D4PHI2X1_L6D4PHI3X2_SP_L5D4PHI2X1_L6D4PHI3X2_wr_en),
.number_out(SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4),
.start(TE_L5D4PHI2X1_L6D4PHI3X2_start),
.done(SP_L5D4PHI2X1_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI3X1_L6D4PHI3X2_SP_L5D4PHI3X1_L6D4PHI3X2;
wire TE_L5D4PHI3X1_L6D4PHI3X2_SP_L5D4PHI3X1_L6D4PHI3X2_wr_en;
wire [5:0] SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3X1_L6D4PHI3X2(
.data_in(TE_L5D4PHI3X1_L6D4PHI3X2_SP_L5D4PHI3X1_L6D4PHI3X2),
.enable(TE_L5D4PHI3X1_L6D4PHI3X2_SP_L5D4PHI3X1_L6D4PHI3X2_wr_en),
.number_out(SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4),
.start(TE_L5D4PHI3X1_L6D4PHI3X2_start),
.done(SP_L5D4PHI3X1_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI3X1_L6D4PHI4X2_SP_L5D4PHI3X1_L6D4PHI4X2;
wire TE_L5D4PHI3X1_L6D4PHI4X2_SP_L5D4PHI3X1_L6D4PHI4X2_wr_en;
wire [5:0] SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3X1_L6D4PHI4X2(
.data_in(TE_L5D4PHI3X1_L6D4PHI4X2_SP_L5D4PHI3X1_L6D4PHI4X2),
.enable(TE_L5D4PHI3X1_L6D4PHI4X2_SP_L5D4PHI3X1_L6D4PHI4X2_wr_en),
.number_out(SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4),
.start(TE_L5D4PHI3X1_L6D4PHI4X2_start),
.done(SP_L5D4PHI3X1_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI1X2_L6D4PHI1X2_SP_L5D4PHI1X2_L6D4PHI1X2;
wire TE_L5D4PHI1X2_L6D4PHI1X2_SP_L5D4PHI1X2_L6D4PHI1X2_wr_en;
wire [5:0] SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1X2_L6D4PHI1X2(
.data_in(TE_L5D4PHI1X2_L6D4PHI1X2_SP_L5D4PHI1X2_L6D4PHI1X2),
.enable(TE_L5D4PHI1X2_L6D4PHI1X2_SP_L5D4PHI1X2_L6D4PHI1X2_wr_en),
.number_out(SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4),
.start(TE_L5D4PHI1X2_L6D4PHI1X2_start),
.done(SP_L5D4PHI1X2_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI1X2_L6D4PHI2X2_SP_L5D4PHI1X2_L6D4PHI2X2;
wire TE_L5D4PHI1X2_L6D4PHI2X2_SP_L5D4PHI1X2_L6D4PHI2X2_wr_en;
wire [5:0] SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI1X2_L6D4PHI2X2(
.data_in(TE_L5D4PHI1X2_L6D4PHI2X2_SP_L5D4PHI1X2_L6D4PHI2X2),
.enable(TE_L5D4PHI1X2_L6D4PHI2X2_SP_L5D4PHI1X2_L6D4PHI2X2_wr_en),
.number_out(SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4),
.start(TE_L5D4PHI1X2_L6D4PHI2X2_start),
.done(SP_L5D4PHI1X2_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI2X2_L6D4PHI2X2_SP_L5D4PHI2X2_L6D4PHI2X2;
wire TE_L5D4PHI2X2_L6D4PHI2X2_SP_L5D4PHI2X2_L6D4PHI2X2_wr_en;
wire [5:0] SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2X2_L6D4PHI2X2(
.data_in(TE_L5D4PHI2X2_L6D4PHI2X2_SP_L5D4PHI2X2_L6D4PHI2X2),
.enable(TE_L5D4PHI2X2_L6D4PHI2X2_SP_L5D4PHI2X2_L6D4PHI2X2_wr_en),
.number_out(SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4),
.start(TE_L5D4PHI2X2_L6D4PHI2X2_start),
.done(SP_L5D4PHI2X2_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI2X2_L6D4PHI3X2_SP_L5D4PHI2X2_L6D4PHI3X2;
wire TE_L5D4PHI2X2_L6D4PHI3X2_SP_L5D4PHI2X2_L6D4PHI3X2_wr_en;
wire [5:0] SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI2X2_L6D4PHI3X2(
.data_in(TE_L5D4PHI2X2_L6D4PHI3X2_SP_L5D4PHI2X2_L6D4PHI3X2),
.enable(TE_L5D4PHI2X2_L6D4PHI3X2_SP_L5D4PHI2X2_L6D4PHI3X2_wr_en),
.number_out(SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4),
.start(TE_L5D4PHI2X2_L6D4PHI3X2_start),
.done(SP_L5D4PHI2X2_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI3X2_L6D4PHI3X2_SP_L5D4PHI3X2_L6D4PHI3X2;
wire TE_L5D4PHI3X2_L6D4PHI3X2_SP_L5D4PHI3X2_L6D4PHI3X2_wr_en;
wire [5:0] SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3X2_L6D4PHI3X2(
.data_in(TE_L5D4PHI3X2_L6D4PHI3X2_SP_L5D4PHI3X2_L6D4PHI3X2),
.enable(TE_L5D4PHI3X2_L6D4PHI3X2_SP_L5D4PHI3X2_L6D4PHI3X2_wr_en),
.number_out(SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4),
.start(TE_L5D4PHI3X2_L6D4PHI3X2_start),
.done(SP_L5D4PHI3X2_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] TE_L5D4PHI3X2_L6D4PHI4X2_SP_L5D4PHI3X2_L6D4PHI4X2;
wire TE_L5D4PHI3X2_L6D4PHI4X2_SP_L5D4PHI3X2_L6D4PHI4X2_wr_en;
wire [5:0] SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4_number;
wire [8:0] SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4_read_add;
wire [11:0] SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4;
StubPairs  SP_L5D4PHI3X2_L6D4PHI4X2(
.data_in(TE_L5D4PHI3X2_L6D4PHI4X2_SP_L5D4PHI3X2_L6D4PHI4X2),
.enable(TE_L5D4PHI3X2_L6D4PHI4X2_SP_L5D4PHI3X2_L6D4PHI4X2_wr_en),
.number_out(SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4_number),
.read_add(SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4_read_add),
.data_out(SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4),
.start(TE_L5D4PHI3X2_L6D4PHI4X2_start),
.done(SP_L5D4PHI3X2_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L5D4_AS_L5D4n1;
wire VMR_L5D4_AS_L5D4n1_wr_en;
wire [10:0] AS_L5D4n1_TC_L5D4L6D4_read_add;
wire [35:0] AS_L5D4n1_TC_L5D4L6D4;
AllStubs  AS_L5D4n1(
.data_in(VMR_L5D4_AS_L5D4n1),
.enable(VMR_L5D4_AS_L5D4n1_wr_en),
.read_add(AS_L5D4n1_TC_L5D4L6D4_read_add),
.data_out(AS_L5D4n1_TC_L5D4L6D4),
.start(VMR_L5D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L6D4_AS_L6D4n2;
wire VMR_L6D4_AS_L6D4n2_wr_en;
wire [10:0] AS_L6D4n2_TC_L5D4L6D4_read_add;
wire [35:0] AS_L6D4n2_TC_L5D4L6D4;
AllStubs  AS_L6D4n2(
.data_in(VMR_L6D4_AS_L6D4n2),
.enable(VMR_L6D4_AS_L6D4n2_wr_en),
.read_add(AS_L6D4n2_TC_L5D4L6D4_read_add),
.data_out(AS_L6D4n2_TC_L5D4L6D4),
.start(VMR_L6D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3;
wire TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D4L6D4_L3(
.data_in(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3),
.enable(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3_wr_en),
.number_out(TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_ToPlus_L5D4L6D4_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3;
wire TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D3L6D4_L3(
.data_in(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3),
.enable(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_ToPlus_L5D3L6D4_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3;
wire TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D3L6D3_L3(
.data_in(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3),
.enable(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_ToPlus_L5D3L6D3_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3;
wire TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L1D4L2D4_L3(
.data_in(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3),
.enable(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3_wr_en),
.number_out(TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus),
.start(TC_L1D4L2D4_proj_start),
.done(TPROJ_ToPlus_L1D4L2D4_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3;
wire TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L1D3L2D4_L3(
.data_in(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3),
.enable(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus),
.start(TC_L1D3L2D4_proj_start),
.done(TPROJ_ToPlus_L1D3L2D4_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3;
wire TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L1D3L2D3_L3(
.data_in(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3),
.enable(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_ToPlus_L1D3L2D3_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4;
wire TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D4L6D4_L4(
.data_in(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4),
.enable(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4_wr_en),
.number_out(TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_ToPlus_L5D4L6D4_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4;
wire TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D3L6D4_L4(
.data_in(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4),
.enable(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_ToPlus_L5D3L6D4_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4;
wire TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D3L6D3_L4(
.data_in(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4),
.enable(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_ToPlus_L5D3L6D3_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4;
wire TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L1D3L2D4_L4(
.data_in(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4),
.enable(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus),
.start(TC_L1D3L2D4_proj_start),
.done(TPROJ_ToPlus_L1D3L2D4_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4;
wire TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L1D3L2D3_L4(
.data_in(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4),
.enable(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_ToPlus_L1D3L2D3_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2;
wire TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D4L6D4_L2(
.data_in(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2),
.enable(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2_wr_en),
.number_out(TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_ToPlus_L5D4L6D4_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2;
wire TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D3L6D4_L2(
.data_in(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2),
.enable(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_ToPlus_L5D3L6D4_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2;
wire TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D3L6D3_L2(
.data_in(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2),
.enable(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_ToPlus_L5D3L6D3_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2;
wire TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D4L4D4_L2(
.data_in(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2),
.enable(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2_wr_en),
.number_out(TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_ToPlus_L3D4L4D4_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2;
wire TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D3L4D4_L2(
.data_in(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2),
.enable(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_ToPlus_L3D3L4D4_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2;
wire TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D3L4D3_L2(
.data_in(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2),
.enable(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_ToPlus_L3D3L4D3_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5;
wire TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D4L4D4_L5(
.data_in(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5),
.enable(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5_wr_en),
.number_out(TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus_number),
.read_add(TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_ToPlus_L3D4L4D4_L5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5;
wire TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D3L4D4_L5(
.data_in(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5),
.enable(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_ToPlus_L3D3L4D4_L5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5;
wire TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D3L4D3_L5(
.data_in(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5),
.enable(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_ToPlus_L3D3L4D3_L5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5;
wire TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L1D3L2D3_L5(
.data_in(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5),
.enable(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_ToPlus_L1D3L2D3_L5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1;
wire TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D4L6D4_L1(
.data_in(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1),
.enable(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1_wr_en),
.number_out(TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_ToPlus_L5D4L6D4_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1;
wire TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D3L6D4_L1(
.data_in(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1),
.enable(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_ToPlus_L5D3L6D4_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1;
wire TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L5D3L6D3_L1(
.data_in(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1),
.enable(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1_wr_en),
.number_out(TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_ToPlus_L5D3L6D3_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1;
wire TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D4L4D4_L1(
.data_in(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1),
.enable(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1_wr_en),
.number_out(TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_ToPlus_L3D4L4D4_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1;
wire TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D3L4D4_L1(
.data_in(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1),
.enable(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_ToPlus_L3D3L4D4_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1;
wire TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D3L4D3_L1(
.data_in(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1),
.enable(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_ToPlus_L3D3L4D3_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6;
wire TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D4L4D4_L6(
.data_in(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6),
.enable(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6_wr_en),
.number_out(TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_ToPlus_L3D4L4D4_L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6;
wire TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D3L4D4_L6(
.data_in(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6),
.enable(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_ToPlus_L3D3L4D4_L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6;
wire TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L3D3L4D3_L6(
.data_in(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6),
.enable(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6_wr_en),
.number_out(TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_ToPlus_L3D3L4D3_L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6;
wire TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6_wr_en;
wire [5:0] TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus_number;
wire [9:0] TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus_read_add;
wire [53:0] TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus;
TrackletProjections #(1'b1) TPROJ_ToPlus_L1D3L2D3_L6(
.data_in(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6),
.enable(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6_wr_en),
.number_out(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus_number),
.read_add(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus_read_add),
.data_out(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_ToPlus_L1D3L2D3_L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3;
wire TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D4L6D4_L3(
.data_in(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3),
.enable(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3_wr_en),
.number_out(TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_ToMinus_L5D4L6D4_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3;
wire TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D3L6D4_L3(
.data_in(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3),
.enable(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_ToMinus_L5D3L6D4_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3;
wire TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D3L6D3_L3(
.data_in(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3),
.enable(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_ToMinus_L5D3L6D3_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3;
wire TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L1D4L2D4_L3(
.data_in(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3),
.enable(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3_wr_en),
.number_out(TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus),
.start(TC_L1D4L2D4_proj_start),
.done(TPROJ_ToMinus_L1D4L2D4_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3;
wire TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L1D3L2D4_L3(
.data_in(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3),
.enable(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus),
.start(TC_L1D3L2D4_proj_start),
.done(TPROJ_ToMinus_L1D3L2D4_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3;
wire TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L1D3L2D3_L3(
.data_in(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3),
.enable(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_ToMinus_L1D3L2D3_L3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4;
wire TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D4L6D4_L4(
.data_in(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4),
.enable(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4_wr_en),
.number_out(TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_ToMinus_L5D4L6D4_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4;
wire TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D3L6D4_L4(
.data_in(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4),
.enable(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_ToMinus_L5D3L6D4_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4;
wire TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D3L6D3_L4(
.data_in(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4),
.enable(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_ToMinus_L5D3L6D3_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4;
wire TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L1D3L2D4_L4(
.data_in(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4),
.enable(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus),
.start(TC_L1D3L2D4_proj_start),
.done(TPROJ_ToMinus_L1D3L2D4_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4;
wire TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L1D3L2D3_L4(
.data_in(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4),
.enable(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_ToMinus_L1D3L2D3_L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2;
wire TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D4L6D4_L2(
.data_in(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2),
.enable(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2_wr_en),
.number_out(TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_ToMinus_L5D4L6D4_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2;
wire TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D3L6D4_L2(
.data_in(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2),
.enable(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_ToMinus_L5D3L6D4_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2;
wire TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D3L6D3_L2(
.data_in(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2),
.enable(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_ToMinus_L5D3L6D3_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2;
wire TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D4L4D4_L2(
.data_in(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2),
.enable(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2_wr_en),
.number_out(TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_ToMinus_L3D4L4D4_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2;
wire TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D3L4D4_L2(
.data_in(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2),
.enable(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_ToMinus_L3D3L4D4_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2;
wire TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D3L4D3_L2(
.data_in(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2),
.enable(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_ToMinus_L3D3L4D3_L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5;
wire TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D4L4D4_L5(
.data_in(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5),
.enable(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5_wr_en),
.number_out(TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus_number),
.read_add(TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_ToMinus_L3D4L4D4_L5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5;
wire TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D3L4D4_L5(
.data_in(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5),
.enable(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_ToMinus_L3D3L4D4_L5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5;
wire TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D3L4D3_L5(
.data_in(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5),
.enable(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_ToMinus_L3D3L4D3_L5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5;
wire TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L1D3L2D3_L5(
.data_in(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5),
.enable(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_ToMinus_L1D3L2D3_L5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1;
wire TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D4L6D4_L1(
.data_in(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1),
.enable(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1_wr_en),
.number_out(TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_ToMinus_L5D4L6D4_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1;
wire TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D3L6D4_L1(
.data_in(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1),
.enable(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_ToMinus_L5D3L6D4_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1;
wire TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L5D3L6D3_L1(
.data_in(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1),
.enable(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1_wr_en),
.number_out(TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_ToMinus_L5D3L6D3_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1;
wire TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D4L4D4_L1(
.data_in(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1),
.enable(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1_wr_en),
.number_out(TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_ToMinus_L3D4L4D4_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1;
wire TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D3L4D4_L1(
.data_in(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1),
.enable(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_ToMinus_L3D3L4D4_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1;
wire TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D3L4D3_L1(
.data_in(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1),
.enable(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_ToMinus_L3D3L4D3_L1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6;
wire TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D4L4D4_L6(
.data_in(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6),
.enable(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6_wr_en),
.number_out(TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_ToMinus_L3D4L4D4_L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6;
wire TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D3L4D4_L6(
.data_in(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6),
.enable(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_ToMinus_L3D3L4D4_L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6;
wire TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L3D3L4D3_L6(
.data_in(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6),
.enable(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6_wr_en),
.number_out(TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_ToMinus_L3D3L4D3_L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6;
wire TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6_wr_en;
wire [5:0] TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus_number;
wire [9:0] TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus_read_add;
wire [53:0] TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus;
TrackletProjections #(1'b1) TPROJ_ToMinus_L1D3L2D3_L6(
.data_in(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6),
.enable(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6_wr_en),
.number_out(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus_number),
.read_add(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus_read_add),
.data_out(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_ToMinus_L1D3L2D3_L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L3L4;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4;
TrackletProjections #(1'b1) TPROJ_FromPlus_L1D3_L3L4(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L3L4),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_number),
.read_add(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_L1D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L3L4;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4;
TrackletProjections #(1'b1) TPROJ_FromMinus_L1D3_L3L4(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L3L4),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_number),
.read_add(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_L1D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L1D3(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3_wr_en),
.number_out(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_L3D3L4D3_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L1D3(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3_wr_en),
.number_out(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_L3D3L4D4_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L1D3(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3_wr_en),
.number_out(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_L3D4L4D4_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L3L4;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4;
TrackletProjections #(1'b1) TPROJ_FromPlus_L2D3_L3L4(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L3L4),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_number),
.read_add(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_L2D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L3L4;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4;
TrackletProjections #(1'b1) TPROJ_FromMinus_L2D3_L3L4(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L3L4),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_number),
.read_add(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_L2D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L2D3(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3_wr_en),
.number_out(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_L3D3L4D3_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L2D3(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3_wr_en),
.number_out(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_L3D3L4D4_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L2D3(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3_wr_en),
.number_out(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_L3D4L4D4_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L3L4;
wire PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_number;
wire [9:0] TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4;
TrackletProjections #(1'b1) TPROJ_FromPlus_L5D3_L3L4(
.data_in(PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L3L4),
.enable(PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_number),
.read_add(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_read_add),
.data_out(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4),
.start(PT_F1L5_Plus_start),
.done(TPROJ_FromPlus_L5D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L3L4;
wire PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_number;
wire [9:0] TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4;
TrackletProjections #(1'b1) TPROJ_FromMinus_L5D3_L3L4(
.data_in(PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L3L4),
.enable(PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_number),
.read_add(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_read_add),
.data_out(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4),
.start(PT_F1L5_Minus_start),
.done(TPROJ_FromMinus_L5D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L5D3(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3_wr_en),
.number_out(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_L3D3L4D3_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L3L4;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_number;
wire [9:0] TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4;
TrackletProjections #(1'b1) TPROJ_FromPlus_L6D3_L3L4(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L3L4),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_number),
.read_add(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_read_add),
.data_out(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_L6D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L3L4;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_number;
wire [9:0] TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4;
TrackletProjections #(1'b1) TPROJ_FromMinus_L6D3_L3L4(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L3L4),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_number),
.read_add(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_read_add),
.data_out(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_L6D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L6D3(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3_wr_en),
.number_out(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_L3D3L4D3_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L3L4;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_number;
wire [9:0] TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4;
TrackletProjections #(1'b1) TPROJ_FromPlus_L1D4_L3L4(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L3L4),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_number),
.read_add(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_read_add),
.data_out(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_L1D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L3L4;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_number;
wire [9:0] TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4;
TrackletProjections #(1'b1) TPROJ_FromMinus_L1D4_L3L4(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L3L4),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_number),
.read_add(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_read_add),
.data_out(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_L1D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L3L4;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_number;
wire [9:0] TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4;
TrackletProjections #(1'b1) TPROJ_FromPlus_L2D4_L3L4(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L3L4),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_number),
.read_add(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_read_add),
.data_out(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_L2D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L3L4;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_number;
wire [9:0] TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4;
TrackletProjections #(1'b1) TPROJ_FromMinus_L2D4_L3L4(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L3L4),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_number),
.read_add(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_read_add),
.data_out(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_L2D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L2D4(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4_wr_en),
.number_out(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_L3D4L4D4_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L3L4;
wire PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4;
TrackletProjections #(1'b1) TPROJ_FromPlus_L5D4_L3L4(
.data_in(PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L3L4),
.enable(PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_number),
.read_add(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4),
.start(PT_F1L5_Plus_start),
.done(TPROJ_FromPlus_L5D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L3L4;
wire PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4;
TrackletProjections #(1'b1) TPROJ_FromMinus_L5D4_L3L4(
.data_in(PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L3L4),
.enable(PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_number),
.read_add(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4),
.start(PT_F1L5_Minus_start),
.done(TPROJ_FromMinus_L5D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L5D4(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4_wr_en),
.number_out(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_L3D3L4D3_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L5D4(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4_wr_en),
.number_out(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_L3D3L4D4_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L5D4(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4_wr_en),
.number_out(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_L3D4L4D4_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L3L4;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L3L4_wr_en;
wire [5:0] TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4;
TrackletProjections #(1'b1) TPROJ_FromPlus_L6D4_L3L4(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L3L4),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L3L4_wr_en),
.number_out(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_number),
.read_add(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_L6D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L3L4;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L3L4_wr_en;
wire [5:0] TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4;
TrackletProjections #(1'b1) TPROJ_FromMinus_L6D4_L3L4(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L3L4),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L3L4_wr_en),
.number_out(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_number),
.read_add(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_L6D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4;
wire TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4_wr_en;
wire [5:0] TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D3_L6D4(
.data_in(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4),
.enable(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4_wr_en),
.number_out(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_number),
.read_add(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4),
.start(TC_L3D3L4D3_proj_start),
.done(TPROJ_L3D3L4D3_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4;
wire TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4_wr_en;
wire [5:0] TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4;
TrackletProjections  TPROJ_L3D3L4D4_L6D4(
.data_in(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4),
.enable(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4_wr_en),
.number_out(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_number),
.read_add(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4),
.start(TC_L3D3L4D4_proj_start),
.done(TPROJ_L3D3L4D4_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4;
wire TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4_wr_en;
wire [5:0] TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_number;
wire [9:0] TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_read_add;
wire [53:0] TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4;
TrackletProjections  TPROJ_L3D4L4D4_L6D4(
.data_in(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4),
.enable(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4_wr_en),
.number_out(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_number),
.read_add(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_read_add),
.data_out(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4),
.start(TC_L3D4L4D4_proj_start),
.done(TPROJ_L3D4L4D4_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L1L2;
wire PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_number;
wire [9:0] TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2;
TrackletProjections #(1'b1) TPROJ_FromPlus_L3D3_L1L2(
.data_in(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L1L2),
.enable(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_number),
.read_add(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_read_add),
.data_out(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2),
.start(PT_L3F3F5_Plus_start),
.done(TPROJ_FromPlus_L3D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L1L2;
wire PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_number;
wire [9:0] TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2;
TrackletProjections #(1'b1) TPROJ_FromMinus_L3D3_L1L2(
.data_in(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L1L2),
.enable(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_number),
.read_add(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_read_add),
.data_out(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2),
.start(PT_L3F3F5_Minus_start),
.done(TPROJ_FromMinus_L3D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L3D3(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3_wr_en),
.number_out(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_L1D3L2D3_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L1L2;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_number;
wire [9:0] TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2;
TrackletProjections #(1'b1) TPROJ_FromPlus_L4D3_L1L2(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L1L2),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_number),
.read_add(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_read_add),
.data_out(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_L4D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L1L2;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_number;
wire [9:0] TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2;
TrackletProjections #(1'b1) TPROJ_FromMinus_L4D3_L1L2(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L1L2),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_number),
.read_add(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_read_add),
.data_out(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_L4D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L4D3(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3_wr_en),
.number_out(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_L1D3L2D3_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L1L2;
wire PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_number;
wire [9:0] TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2;
TrackletProjections #(1'b1) TPROJ_FromPlus_L5D3_L1L2(
.data_in(PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L1L2),
.enable(PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_number),
.read_add(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_read_add),
.data_out(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2),
.start(PT_F1L5_Plus_start),
.done(TPROJ_FromPlus_L5D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L1L2;
wire PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_number;
wire [9:0] TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2;
TrackletProjections #(1'b1) TPROJ_FromMinus_L5D3_L1L2(
.data_in(PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L1L2),
.enable(PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_number),
.read_add(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_read_add),
.data_out(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2),
.start(PT_F1L5_Minus_start),
.done(TPROJ_FromMinus_L5D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L5D3(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3_wr_en),
.number_out(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_L1D3L2D3_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L1L2;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_number;
wire [9:0] TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2;
TrackletProjections #(1'b1) TPROJ_FromPlus_L6D3_L1L2(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L1L2),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_number),
.read_add(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_read_add),
.data_out(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_L6D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L1L2;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_number;
wire [9:0] TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2;
TrackletProjections #(1'b1) TPROJ_FromMinus_L6D3_L1L2(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L1L2),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_number),
.read_add(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_read_add),
.data_out(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_L6D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L6D3(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3_wr_en),
.number_out(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_L1D3L2D3_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L1L2;
wire PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2;
TrackletProjections #(1'b1) TPROJ_FromPlus_L3D4_L1L2(
.data_in(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L1L2),
.enable(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_number),
.read_add(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2),
.start(PT_L3F3F5_Plus_start),
.done(TPROJ_FromPlus_L3D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L1L2;
wire PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2;
TrackletProjections #(1'b1) TPROJ_FromMinus_L3D4_L1L2(
.data_in(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L1L2),
.enable(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_number),
.read_add(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2),
.start(PT_L3F3F5_Minus_start),
.done(TPROJ_FromMinus_L3D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L3D4(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4_wr_en),
.number_out(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_L1D3L2D3_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L3D4(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4_wr_en),
.number_out(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2),
.start(TC_L1D3L2D4_proj_start),
.done(TPROJ_L1D3L2D4_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4;
wire TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4_wr_en;
wire [5:0] TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_number;
wire [9:0] TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_read_add;
wire [53:0] TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2;
TrackletProjections  TPROJ_L1D4L2D4_L3D4(
.data_in(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4),
.enable(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4_wr_en),
.number_out(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_number),
.read_add(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_read_add),
.data_out(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2),
.start(TC_L1D4L2D4_proj_start),
.done(TPROJ_L1D4L2D4_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L1L2;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2;
TrackletProjections #(1'b1) TPROJ_FromPlus_L4D4_L1L2(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L1L2),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_number),
.read_add(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_L4D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L1L2;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2;
TrackletProjections #(1'b1) TPROJ_FromMinus_L4D4_L1L2(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L1L2),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_number),
.read_add(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_L4D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L4D4(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4_wr_en),
.number_out(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_L1D3L2D3_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4;
wire TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4_wr_en;
wire [5:0] TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D4_L4D4(
.data_in(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4),
.enable(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4_wr_en),
.number_out(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_number),
.read_add(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2),
.start(TC_L1D3L2D4_proj_start),
.done(TPROJ_L1D3L2D4_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L1L2;
wire PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_number;
wire [9:0] TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2;
TrackletProjections #(1'b1) TPROJ_FromPlus_L5D4_L1L2(
.data_in(PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L1L2),
.enable(PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_number),
.read_add(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_read_add),
.data_out(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2),
.start(PT_F1L5_Plus_start),
.done(TPROJ_FromPlus_L5D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L1L2;
wire PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_number;
wire [9:0] TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2;
TrackletProjections #(1'b1) TPROJ_FromMinus_L5D4_L1L2(
.data_in(PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L1L2),
.enable(PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_number),
.read_add(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_read_add),
.data_out(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2),
.start(PT_F1L5_Minus_start),
.done(TPROJ_FromMinus_L5D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L5D4(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4_wr_en),
.number_out(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_L1D3L2D3_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L1L2;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L1L2_wr_en;
wire [5:0] TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_number;
wire [9:0] TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_read_add;
wire [53:0] TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2;
TrackletProjections #(1'b1) TPROJ_FromPlus_L6D4_L1L2(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L1L2),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L1L2_wr_en),
.number_out(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_number),
.read_add(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_read_add),
.data_out(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_L6D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L1L2;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L1L2_wr_en;
wire [5:0] TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_number;
wire [9:0] TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_read_add;
wire [53:0] TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2;
TrackletProjections #(1'b1) TPROJ_FromMinus_L6D4_L1L2(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L1L2),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L1L2_wr_en),
.number_out(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_number),
.read_add(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_read_add),
.data_out(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_L6D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4;
wire TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4_wr_en;
wire [5:0] TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_number;
wire [9:0] TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_read_add;
wire [53:0] TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2;
TrackletProjections  TPROJ_L1D3L2D3_L6D4(
.data_in(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4),
.enable(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4_wr_en),
.number_out(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_number),
.read_add(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_read_add),
.data_out(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2),
.start(TC_L1D3L2D3_proj_start),
.done(TPROJ_L1D3L2D3_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L5L6;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6;
TrackletProjections #(1'b1) TPROJ_FromPlus_L1D3_L5L6(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L5L6),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_number),
.read_add(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_L1D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L5L6;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6;
TrackletProjections #(1'b1) TPROJ_FromMinus_L1D3_L5L6(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L5L6),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_number),
.read_add(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_L1D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L1D3(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3_wr_en),
.number_out(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_L5D3L6D3_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L1D3(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3_wr_en),
.number_out(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_L5D3L6D4_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L1D3(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3_wr_en),
.number_out(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_L5D4L6D4_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L5L6;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6;
TrackletProjections #(1'b1) TPROJ_FromPlus_L2D3_L5L6(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L5L6),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_number),
.read_add(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_L2D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L5L6;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6;
TrackletProjections #(1'b1) TPROJ_FromMinus_L2D3_L5L6(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L5L6),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_number),
.read_add(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_L2D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L2D3(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3_wr_en),
.number_out(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_L5D3L6D3_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L2D3(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3_wr_en),
.number_out(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_L5D3L6D4_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L2D3(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3_wr_en),
.number_out(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_L5D4L6D4_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L5L6;
wire PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6;
TrackletProjections #(1'b1) TPROJ_FromPlus_L3D3_L5L6(
.data_in(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L5L6),
.enable(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_number),
.read_add(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6),
.start(PT_L3F3F5_Plus_start),
.done(TPROJ_FromPlus_L3D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L5L6;
wire PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6;
TrackletProjections #(1'b1) TPROJ_FromMinus_L3D3_L5L6(
.data_in(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L5L6),
.enable(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_number),
.read_add(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6),
.start(PT_L3F3F5_Minus_start),
.done(TPROJ_FromMinus_L3D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L3D3(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3_wr_en),
.number_out(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_L5D3L6D3_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L3D3(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3_wr_en),
.number_out(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_L5D3L6D4_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L3D3(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3_wr_en),
.number_out(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_L5D4L6D4_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L5L6;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6;
TrackletProjections #(1'b1) TPROJ_FromPlus_L4D3_L5L6(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L5L6),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_number),
.read_add(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_L4D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L5L6;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6;
TrackletProjections #(1'b1) TPROJ_FromMinus_L4D3_L5L6(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L5L6),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_number),
.read_add(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_L4D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3;
wire TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3_wr_en;
wire [5:0] TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D3_L4D3(
.data_in(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3),
.enable(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3_wr_en),
.number_out(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_number),
.read_add(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6),
.start(TC_L5D3L6D3_proj_start),
.done(TPROJ_L5D3L6D3_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3;
wire TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3_wr_en;
wire [5:0] TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6;
TrackletProjections  TPROJ_L5D3L6D4_L4D3(
.data_in(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3),
.enable(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3_wr_en),
.number_out(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_number),
.read_add(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6),
.start(TC_L5D3L6D4_proj_start),
.done(TPROJ_L5D3L6D4_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L4D3(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3_wr_en),
.number_out(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_L5D4L6D4_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L5L6;
wire PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_number;
wire [9:0] TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6;
TrackletProjections #(1'b1) TPROJ_FromPlus_L1D4_L5L6(
.data_in(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L5L6),
.enable(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_number),
.read_add(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_read_add),
.data_out(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6),
.start(PT_L1L6F4_Plus_start),
.done(TPROJ_FromPlus_L1D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L5L6;
wire PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_number;
wire [9:0] TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6;
TrackletProjections #(1'b1) TPROJ_FromMinus_L1D4_L5L6(
.data_in(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L5L6),
.enable(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_number),
.read_add(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_read_add),
.data_out(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6),
.start(PT_L1L6F4_Minus_start),
.done(TPROJ_FromMinus_L1D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L5L6;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_number;
wire [9:0] TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6;
TrackletProjections #(1'b1) TPROJ_FromPlus_L2D4_L5L6(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L5L6),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_number),
.read_add(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_read_add),
.data_out(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_L2D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L5L6;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_number;
wire [9:0] TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6;
TrackletProjections #(1'b1) TPROJ_FromMinus_L2D4_L5L6(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L5L6),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_number),
.read_add(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_read_add),
.data_out(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_L2D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L5L6;
wire PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_number;
wire [9:0] TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6;
TrackletProjections #(1'b1) TPROJ_FromPlus_L3D4_L5L6(
.data_in(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L5L6),
.enable(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_number),
.read_add(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_read_add),
.data_out(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6),
.start(PT_L3F3F5_Plus_start),
.done(TPROJ_FromPlus_L3D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L5L6;
wire PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_number;
wire [9:0] TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6;
TrackletProjections #(1'b1) TPROJ_FromMinus_L3D4_L5L6(
.data_in(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L5L6),
.enable(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_number),
.read_add(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_read_add),
.data_out(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6),
.start(PT_L3F3F5_Minus_start),
.done(TPROJ_FromMinus_L3D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L3D4(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4_wr_en),
.number_out(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_L5D4L6D4_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L5L6;
wire PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L5L6_wr_en;
wire [5:0] TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_number;
wire [9:0] TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_read_add;
wire [53:0] TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6;
TrackletProjections #(1'b1) TPROJ_FromPlus_L4D4_L5L6(
.data_in(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L5L6),
.enable(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L5L6_wr_en),
.number_out(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_number),
.read_add(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_read_add),
.data_out(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6),
.start(PT_L2L4F2_Plus_start),
.done(TPROJ_FromPlus_L4D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L5L6;
wire PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L5L6_wr_en;
wire [5:0] TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_number;
wire [9:0] TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_read_add;
wire [53:0] TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6;
TrackletProjections #(1'b1) TPROJ_FromMinus_L4D4_L5L6(
.data_in(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L5L6),
.enable(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L5L6_wr_en),
.number_out(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_number),
.read_add(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_read_add),
.data_out(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6),
.start(PT_L2L4F2_Minus_start),
.done(TPROJ_FromMinus_L4D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [53:0] TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4;
wire TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4_wr_en;
wire [5:0] TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_number;
wire [9:0] TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_read_add;
wire [53:0] TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6;
TrackletProjections  TPROJ_L5D4L6D4_L4D4(
.data_in(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4),
.enable(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4_wr_en),
.number_out(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_number),
.read_add(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_read_add),
.data_out(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6),
.start(TC_L5D4L6D4_proj_start),
.done(TPROJ_L5D4L6D4_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X1;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1_read_add;
wire [13:0] VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1;
VMProjections  VMPROJ_L3L4_L1D3PHI1X1(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X1),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X1_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1_number),
.read_add(VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1),
.start(PR_L1D3_L3L4_start),
.done(VMPROJ_L3L4_L1D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X1n7;
wire VMR_L1D3_VMS_L1D3PHI1X1n7_wr_en;
wire [5:0] VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1_number;
wire [10:0] VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1_read_add;
wire [18:0] VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1;
VMStubs #("Match") VMS_L1D3PHI1X1n7(
.data_in(VMR_L1D3_VMS_L1D3PHI1X1n7),
.enable(VMR_L1D3_VMS_L1D3PHI1X1n7_wr_en),
.number_out(VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1_number),
.read_add(VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1_read_add),
.data_out(VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X1n7_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X2;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2_read_add;
wire [13:0] VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2;
VMProjections  VMPROJ_L3L4_L1D3PHI1X2(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X2),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X2_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2_number),
.read_add(VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2),
.start(PR_L1D3_L3L4_start),
.done(VMPROJ_L3L4_L1D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X2n7;
wire VMR_L1D3_VMS_L1D3PHI1X2n7_wr_en;
wire [5:0] VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2_number;
wire [10:0] VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2_read_add;
wire [18:0] VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2;
VMStubs #("Match") VMS_L1D3PHI1X2n7(
.data_in(VMR_L1D3_VMS_L1D3PHI1X2n7),
.enable(VMR_L1D3_VMS_L1D3PHI1X2n7_wr_en),
.number_out(VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2_number),
.read_add(VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2_read_add),
.data_out(VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X2n7_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X1;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1_read_add;
wire [13:0] VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1;
VMProjections  VMPROJ_L3L4_L1D3PHI2X1(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X1),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X1_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1_number),
.read_add(VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1),
.start(PR_L1D3_L3L4_start),
.done(VMPROJ_L3L4_L1D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X1n7;
wire VMR_L1D3_VMS_L1D3PHI2X1n7_wr_en;
wire [5:0] VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1_number;
wire [10:0] VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1_read_add;
wire [18:0] VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1;
VMStubs #("Match") VMS_L1D3PHI2X1n7(
.data_in(VMR_L1D3_VMS_L1D3PHI2X1n7),
.enable(VMR_L1D3_VMS_L1D3PHI2X1n7_wr_en),
.number_out(VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1_number),
.read_add(VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1_read_add),
.data_out(VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X1n7_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X2;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2_read_add;
wire [13:0] VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2;
VMProjections  VMPROJ_L3L4_L1D3PHI2X2(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X2),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X2_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2_number),
.read_add(VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2),
.start(PR_L1D3_L3L4_start),
.done(VMPROJ_L3L4_L1D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X2n7;
wire VMR_L1D3_VMS_L1D3PHI2X2n7_wr_en;
wire [5:0] VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2_number;
wire [10:0] VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2_read_add;
wire [18:0] VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2;
VMStubs #("Match") VMS_L1D3PHI2X2n7(
.data_in(VMR_L1D3_VMS_L1D3PHI2X2n7),
.enable(VMR_L1D3_VMS_L1D3PHI2X2n7_wr_en),
.number_out(VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2_number),
.read_add(VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2_read_add),
.data_out(VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X2n7_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X1;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1_read_add;
wire [13:0] VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1;
VMProjections  VMPROJ_L3L4_L1D3PHI3X1(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X1),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X1_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1_number),
.read_add(VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1),
.start(PR_L1D3_L3L4_start),
.done(VMPROJ_L3L4_L1D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X1n7;
wire VMR_L1D3_VMS_L1D3PHI3X1n7_wr_en;
wire [5:0] VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1_number;
wire [10:0] VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1_read_add;
wire [18:0] VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1;
VMStubs #("Match") VMS_L1D3PHI3X1n7(
.data_in(VMR_L1D3_VMS_L1D3PHI3X1n7),
.enable(VMR_L1D3_VMS_L1D3PHI3X1n7_wr_en),
.number_out(VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1_number),
.read_add(VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1_read_add),
.data_out(VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X1n7_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X2;
wire PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2_number;
wire [8:0] VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2_read_add;
wire [13:0] VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2;
VMProjections  VMPROJ_L3L4_L1D3PHI3X2(
.data_in(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X2),
.enable(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X2_wr_en),
.number_out(VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2_number),
.read_add(VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2_read_add),
.data_out(VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2),
.start(PR_L1D3_L3L4_start),
.done(VMPROJ_L3L4_L1D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X2n7;
wire VMR_L1D3_VMS_L1D3PHI3X2n7_wr_en;
wire [5:0] VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2_number;
wire [10:0] VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2_read_add;
wire [18:0] VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2;
VMStubs #("Match") VMS_L1D3PHI3X2n7(
.data_in(VMR_L1D3_VMS_L1D3PHI3X2n7),
.enable(VMR_L1D3_VMS_L1D3PHI3X2n7_wr_en),
.number_out(VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2_number),
.read_add(VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2_read_add),
.data_out(VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X2n7_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X1;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1_read_add;
wire [13:0] VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1;
VMProjections  VMPROJ_L3L4_L1D4PHI1X1(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X1),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X1_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1_number),
.read_add(VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1),
.start(PR_L1D4_L3L4_start),
.done(VMPROJ_L3L4_L1D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI1X1n3;
wire VMR_L1D4_VMS_L1D4PHI1X1n3_wr_en;
wire [5:0] VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1_number;
wire [10:0] VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1_read_add;
wire [18:0] VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1;
VMStubs #("Match") VMS_L1D4PHI1X1n3(
.data_in(VMR_L1D4_VMS_L1D4PHI1X1n3),
.enable(VMR_L1D4_VMS_L1D4PHI1X1n3_wr_en),
.number_out(VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1_number),
.read_add(VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1_read_add),
.data_out(VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X2;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2_read_add;
wire [13:0] VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2;
VMProjections  VMPROJ_L3L4_L1D4PHI1X2(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X2),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X2_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2_number),
.read_add(VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2),
.start(PR_L1D4_L3L4_start),
.done(VMPROJ_L3L4_L1D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI1X2n1;
wire VMR_L1D4_VMS_L1D4PHI1X2n1_wr_en;
wire [5:0] VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2_number;
wire [10:0] VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2_read_add;
wire [18:0] VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2;
VMStubs #("Match") VMS_L1D4PHI1X2n1(
.data_in(VMR_L1D4_VMS_L1D4PHI1X2n1),
.enable(VMR_L1D4_VMS_L1D4PHI1X2n1_wr_en),
.number_out(VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2_number),
.read_add(VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2_read_add),
.data_out(VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI1X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X1;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1_read_add;
wire [13:0] VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1;
VMProjections  VMPROJ_L3L4_L1D4PHI2X1(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X1),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X1_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1_number),
.read_add(VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1),
.start(PR_L1D4_L3L4_start),
.done(VMPROJ_L3L4_L1D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI2X1n3;
wire VMR_L1D4_VMS_L1D4PHI2X1n3_wr_en;
wire [5:0] VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1_number;
wire [10:0] VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1_read_add;
wire [18:0] VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1;
VMStubs #("Match") VMS_L1D4PHI2X1n3(
.data_in(VMR_L1D4_VMS_L1D4PHI2X1n3),
.enable(VMR_L1D4_VMS_L1D4PHI2X1n3_wr_en),
.number_out(VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1_number),
.read_add(VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1_read_add),
.data_out(VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X2;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2_read_add;
wire [13:0] VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2;
VMProjections  VMPROJ_L3L4_L1D4PHI2X2(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X2),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X2_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2_number),
.read_add(VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2),
.start(PR_L1D4_L3L4_start),
.done(VMPROJ_L3L4_L1D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI2X2n1;
wire VMR_L1D4_VMS_L1D4PHI2X2n1_wr_en;
wire [5:0] VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2_number;
wire [10:0] VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2_read_add;
wire [18:0] VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2;
VMStubs #("Match") VMS_L1D4PHI2X2n1(
.data_in(VMR_L1D4_VMS_L1D4PHI2X2n1),
.enable(VMR_L1D4_VMS_L1D4PHI2X2n1_wr_en),
.number_out(VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2_number),
.read_add(VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2_read_add),
.data_out(VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI2X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X1;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1_read_add;
wire [13:0] VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1;
VMProjections  VMPROJ_L3L4_L1D4PHI3X1(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X1),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X1_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1_number),
.read_add(VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1),
.start(PR_L1D4_L3L4_start),
.done(VMPROJ_L3L4_L1D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI3X1n3;
wire VMR_L1D4_VMS_L1D4PHI3X1n3_wr_en;
wire [5:0] VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1_number;
wire [10:0] VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1_read_add;
wire [18:0] VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1;
VMStubs #("Match") VMS_L1D4PHI3X1n3(
.data_in(VMR_L1D4_VMS_L1D4PHI3X1n3),
.enable(VMR_L1D4_VMS_L1D4PHI3X1n3_wr_en),
.number_out(VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1_number),
.read_add(VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1_read_add),
.data_out(VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X2;
wire PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2_number;
wire [8:0] VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2_read_add;
wire [13:0] VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2;
VMProjections  VMPROJ_L3L4_L1D4PHI3X2(
.data_in(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X2),
.enable(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X2_wr_en),
.number_out(VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2_number),
.read_add(VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2_read_add),
.data_out(VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2),
.start(PR_L1D4_L3L4_start),
.done(VMPROJ_L3L4_L1D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI3X2n1;
wire VMR_L1D4_VMS_L1D4PHI3X2n1_wr_en;
wire [5:0] VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2_number;
wire [10:0] VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2_read_add;
wire [18:0] VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2;
VMStubs #("Match") VMS_L1D4PHI3X2n1(
.data_in(VMR_L1D4_VMS_L1D4PHI3X2n1),
.enable(VMR_L1D4_VMS_L1D4PHI3X2n1_wr_en),
.number_out(VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2_number),
.read_add(VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2_read_add),
.data_out(VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI3X2n1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X1;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1_read_add;
wire [13:0] VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1;
VMProjections  VMPROJ_L3L4_L2D3PHI1X1(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X1),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X1_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1_number),
.read_add(VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1),
.start(PR_L2D3_L3L4_start),
.done(VMPROJ_L3L4_L2D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI1X1n2;
wire VMR_L2D3_VMS_L2D3PHI1X1n2_wr_en;
wire [5:0] VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1_number;
wire [10:0] VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1_read_add;
wire [18:0] VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1;
VMStubs #("Match") VMS_L2D3PHI1X1n2(
.data_in(VMR_L2D3_VMS_L2D3PHI1X1n2),
.enable(VMR_L2D3_VMS_L2D3PHI1X1n2_wr_en),
.number_out(VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1_number),
.read_add(VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1_read_add),
.data_out(VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X2;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2_read_add;
wire [13:0] VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2;
VMProjections  VMPROJ_L3L4_L2D3PHI1X2(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X2),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X2_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2_number),
.read_add(VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2),
.start(PR_L2D3_L3L4_start),
.done(VMPROJ_L3L4_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI1X2n3;
wire VMR_L2D3_VMS_L2D3PHI1X2n3_wr_en;
wire [5:0] VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2_number;
wire [10:0] VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2_read_add;
wire [18:0] VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2;
VMStubs #("Match") VMS_L2D3PHI1X2n3(
.data_in(VMR_L2D3_VMS_L2D3PHI1X2n3),
.enable(VMR_L2D3_VMS_L2D3PHI1X2n3_wr_en),
.number_out(VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2_number),
.read_add(VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2_read_add),
.data_out(VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X1;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1_read_add;
wire [13:0] VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1;
VMProjections  VMPROJ_L3L4_L2D3PHI2X1(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X1),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X1_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1_number),
.read_add(VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1),
.start(PR_L2D3_L3L4_start),
.done(VMPROJ_L3L4_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X1n3;
wire VMR_L2D3_VMS_L2D3PHI2X1n3_wr_en;
wire [5:0] VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1_number;
wire [10:0] VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1_read_add;
wire [18:0] VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1;
VMStubs #("Match") VMS_L2D3PHI2X1n3(
.data_in(VMR_L2D3_VMS_L2D3PHI2X1n3),
.enable(VMR_L2D3_VMS_L2D3PHI2X1n3_wr_en),
.number_out(VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1_number),
.read_add(VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1_read_add),
.data_out(VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X2;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2_read_add;
wire [13:0] VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2;
VMProjections  VMPROJ_L3L4_L2D3PHI2X2(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X2),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X2_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2_number),
.read_add(VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2),
.start(PR_L2D3_L3L4_start),
.done(VMPROJ_L3L4_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X2n5;
wire VMR_L2D3_VMS_L2D3PHI2X2n5_wr_en;
wire [5:0] VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2_number;
wire [10:0] VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2_read_add;
wire [18:0] VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2;
VMStubs #("Match") VMS_L2D3PHI2X2n5(
.data_in(VMR_L2D3_VMS_L2D3PHI2X2n5),
.enable(VMR_L2D3_VMS_L2D3PHI2X2n5_wr_en),
.number_out(VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2_number),
.read_add(VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2_read_add),
.data_out(VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X1;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1_read_add;
wire [13:0] VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1;
VMProjections  VMPROJ_L3L4_L2D3PHI3X1(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X1),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X1_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1_number),
.read_add(VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1),
.start(PR_L2D3_L3L4_start),
.done(VMPROJ_L3L4_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X1n3;
wire VMR_L2D3_VMS_L2D3PHI3X1n3_wr_en;
wire [5:0] VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1_number;
wire [10:0] VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1_read_add;
wire [18:0] VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1;
VMStubs #("Match") VMS_L2D3PHI3X1n3(
.data_in(VMR_L2D3_VMS_L2D3PHI3X1n3),
.enable(VMR_L2D3_VMS_L2D3PHI3X1n3_wr_en),
.number_out(VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1_number),
.read_add(VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1_read_add),
.data_out(VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X2;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2_read_add;
wire [13:0] VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2;
VMProjections  VMPROJ_L3L4_L2D3PHI3X2(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X2),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X2_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2_number),
.read_add(VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2),
.start(PR_L2D3_L3L4_start),
.done(VMPROJ_L3L4_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X2n5;
wire VMR_L2D3_VMS_L2D3PHI3X2n5_wr_en;
wire [5:0] VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2_number;
wire [10:0] VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2_read_add;
wire [18:0] VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2;
VMStubs #("Match") VMS_L2D3PHI3X2n5(
.data_in(VMR_L2D3_VMS_L2D3PHI3X2n5),
.enable(VMR_L2D3_VMS_L2D3PHI3X2n5_wr_en),
.number_out(VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2_number),
.read_add(VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2_read_add),
.data_out(VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X1;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1_read_add;
wire [13:0] VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1;
VMProjections  VMPROJ_L3L4_L2D3PHI4X1(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X1),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X1_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1_number),
.read_add(VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1),
.start(PR_L2D3_L3L4_start),
.done(VMPROJ_L3L4_L2D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI4X1n2;
wire VMR_L2D3_VMS_L2D3PHI4X1n2_wr_en;
wire [5:0] VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1_number;
wire [10:0] VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1_read_add;
wire [18:0] VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1;
VMStubs #("Match") VMS_L2D3PHI4X1n2(
.data_in(VMR_L2D3_VMS_L2D3PHI4X1n2),
.enable(VMR_L2D3_VMS_L2D3PHI4X1n2_wr_en),
.number_out(VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1_number),
.read_add(VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1_read_add),
.data_out(VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X2;
wire PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2_number;
wire [8:0] VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2_read_add;
wire [13:0] VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2;
VMProjections  VMPROJ_L3L4_L2D3PHI4X2(
.data_in(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X2),
.enable(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X2_wr_en),
.number_out(VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2_number),
.read_add(VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2_read_add),
.data_out(VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2),
.start(PR_L2D3_L3L4_start),
.done(VMPROJ_L3L4_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI4X2n3;
wire VMR_L2D3_VMS_L2D3PHI4X2n3_wr_en;
wire [5:0] VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2_number;
wire [10:0] VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2_read_add;
wire [18:0] VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2;
VMStubs #("Match") VMS_L2D3PHI4X2n3(
.data_in(VMR_L2D3_VMS_L2D3PHI4X2n3),
.enable(VMR_L2D3_VMS_L2D3PHI4X2n3_wr_en),
.number_out(VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2_number),
.read_add(VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2_read_add),
.data_out(VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI4X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X1;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1_read_add;
wire [13:0] VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1;
VMProjections  VMPROJ_L3L4_L2D4PHI1X1(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X1),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X1_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1_number),
.read_add(VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1),
.start(PR_L2D4_L3L4_start),
.done(VMPROJ_L3L4_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI1X1n3;
wire VMR_L2D4_VMS_L2D4PHI1X1n3_wr_en;
wire [5:0] VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1_number;
wire [10:0] VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1_read_add;
wire [18:0] VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1;
VMStubs #("Match") VMS_L2D4PHI1X1n3(
.data_in(VMR_L2D4_VMS_L2D4PHI1X1n3),
.enable(VMR_L2D4_VMS_L2D4PHI1X1n3_wr_en),
.number_out(VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1_number),
.read_add(VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1_read_add),
.data_out(VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X2;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2_read_add;
wire [13:0] VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2;
VMProjections  VMPROJ_L3L4_L2D4PHI1X2(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X2),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X2_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2_number),
.read_add(VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2),
.start(PR_L2D4_L3L4_start),
.done(VMPROJ_L3L4_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI1X2n3;
wire VMR_L2D4_VMS_L2D4PHI1X2n3_wr_en;
wire [5:0] VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2_number;
wire [10:0] VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2_read_add;
wire [18:0] VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2;
VMStubs #("Match") VMS_L2D4PHI1X2n3(
.data_in(VMR_L2D4_VMS_L2D4PHI1X2n3),
.enable(VMR_L2D4_VMS_L2D4PHI1X2n3_wr_en),
.number_out(VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2_number),
.read_add(VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2_read_add),
.data_out(VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X1;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1_read_add;
wire [13:0] VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1;
VMProjections  VMPROJ_L3L4_L2D4PHI2X1(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X1),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X1_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1_number),
.read_add(VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1),
.start(PR_L2D4_L3L4_start),
.done(VMPROJ_L3L4_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X1n5;
wire VMR_L2D4_VMS_L2D4PHI2X1n5_wr_en;
wire [5:0] VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1_number;
wire [10:0] VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1_read_add;
wire [18:0] VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1;
VMStubs #("Match") VMS_L2D4PHI2X1n5(
.data_in(VMR_L2D4_VMS_L2D4PHI2X1n5),
.enable(VMR_L2D4_VMS_L2D4PHI2X1n5_wr_en),
.number_out(VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1_number),
.read_add(VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1_read_add),
.data_out(VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X2;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2_read_add;
wire [13:0] VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2;
VMProjections  VMPROJ_L3L4_L2D4PHI2X2(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X2),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X2_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2_number),
.read_add(VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2),
.start(PR_L2D4_L3L4_start),
.done(VMPROJ_L3L4_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X2n5;
wire VMR_L2D4_VMS_L2D4PHI2X2n5_wr_en;
wire [5:0] VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2_number;
wire [10:0] VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2_read_add;
wire [18:0] VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2;
VMStubs #("Match") VMS_L2D4PHI2X2n5(
.data_in(VMR_L2D4_VMS_L2D4PHI2X2n5),
.enable(VMR_L2D4_VMS_L2D4PHI2X2n5_wr_en),
.number_out(VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2_number),
.read_add(VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2_read_add),
.data_out(VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X1;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1_read_add;
wire [13:0] VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1;
VMProjections  VMPROJ_L3L4_L2D4PHI3X1(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X1),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X1_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1_number),
.read_add(VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1),
.start(PR_L2D4_L3L4_start),
.done(VMPROJ_L3L4_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X1n5;
wire VMR_L2D4_VMS_L2D4PHI3X1n5_wr_en;
wire [5:0] VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1_number;
wire [10:0] VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1_read_add;
wire [18:0] VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1;
VMStubs #("Match") VMS_L2D4PHI3X1n5(
.data_in(VMR_L2D4_VMS_L2D4PHI3X1n5),
.enable(VMR_L2D4_VMS_L2D4PHI3X1n5_wr_en),
.number_out(VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1_number),
.read_add(VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1_read_add),
.data_out(VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X2;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2_read_add;
wire [13:0] VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2;
VMProjections  VMPROJ_L3L4_L2D4PHI3X2(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X2),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X2_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2_number),
.read_add(VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2),
.start(PR_L2D4_L3L4_start),
.done(VMPROJ_L3L4_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X2n5;
wire VMR_L2D4_VMS_L2D4PHI3X2n5_wr_en;
wire [5:0] VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2_number;
wire [10:0] VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2_read_add;
wire [18:0] VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2;
VMStubs #("Match") VMS_L2D4PHI3X2n5(
.data_in(VMR_L2D4_VMS_L2D4PHI3X2n5),
.enable(VMR_L2D4_VMS_L2D4PHI3X2n5_wr_en),
.number_out(VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2_number),
.read_add(VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2_read_add),
.data_out(VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X1;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X1_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1_read_add;
wire [13:0] VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1;
VMProjections  VMPROJ_L3L4_L2D4PHI4X1(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X1),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X1_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1_number),
.read_add(VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1),
.start(PR_L2D4_L3L4_start),
.done(VMPROJ_L3L4_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI4X1n3;
wire VMR_L2D4_VMS_L2D4PHI4X1n3_wr_en;
wire [5:0] VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1_number;
wire [10:0] VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1_read_add;
wire [18:0] VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1;
VMStubs #("Match") VMS_L2D4PHI4X1n3(
.data_in(VMR_L2D4_VMS_L2D4PHI4X1n3),
.enable(VMR_L2D4_VMS_L2D4PHI4X1n3_wr_en),
.number_out(VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1_number),
.read_add(VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1_read_add),
.data_out(VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI4X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X2;
wire PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X2_wr_en;
wire [5:0] VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2_number;
wire [8:0] VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2_read_add;
wire [13:0] VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2;
VMProjections  VMPROJ_L3L4_L2D4PHI4X2(
.data_in(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X2),
.enable(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X2_wr_en),
.number_out(VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2_number),
.read_add(VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2_read_add),
.data_out(VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2),
.start(PR_L2D4_L3L4_start),
.done(VMPROJ_L3L4_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI4X2n3;
wire VMR_L2D4_VMS_L2D4PHI4X2n3_wr_en;
wire [5:0] VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2_number;
wire [10:0] VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2_read_add;
wire [18:0] VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2;
VMStubs #("Match") VMS_L2D4PHI4X2n3(
.data_in(VMR_L2D4_VMS_L2D4PHI4X2n3),
.enable(VMR_L2D4_VMS_L2D4PHI4X2n3_wr_en),
.number_out(VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2_number),
.read_add(VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2_read_add),
.data_out(VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI4X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X1;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1_read_add;
wire [13:0] VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1;
VMProjections  VMPROJ_L3L4_L5D3PHI1X1(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X1),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X1_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1_number),
.read_add(VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1),
.start(PR_L5D3_L3L4_start),
.done(VMPROJ_L3L4_L5D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X1n5;
wire VMR_L5D3_VMS_L5D3PHI1X1n5_wr_en;
wire [5:0] VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1_number;
wire [10:0] VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1_read_add;
wire [18:0] VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1;
VMStubs #("Match") VMS_L5D3PHI1X1n5(
.data_in(VMR_L5D3_VMS_L5D3PHI1X1n5),
.enable(VMR_L5D3_VMS_L5D3PHI1X1n5_wr_en),
.number_out(VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1_number),
.read_add(VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1_read_add),
.data_out(VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X2;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2_read_add;
wire [13:0] VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2;
VMProjections  VMPROJ_L3L4_L5D3PHI1X2(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X2),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X2_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2_number),
.read_add(VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2),
.start(PR_L5D3_L3L4_start),
.done(VMPROJ_L3L4_L5D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X2n5;
wire VMR_L5D3_VMS_L5D3PHI1X2n5_wr_en;
wire [5:0] VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2_number;
wire [10:0] VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2_read_add;
wire [18:0] VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2;
VMStubs #("Match") VMS_L5D3PHI1X2n5(
.data_in(VMR_L5D3_VMS_L5D3PHI1X2n5),
.enable(VMR_L5D3_VMS_L5D3PHI1X2n5_wr_en),
.number_out(VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2_number),
.read_add(VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2_read_add),
.data_out(VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X1;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1_read_add;
wire [13:0] VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1;
VMProjections  VMPROJ_L3L4_L5D3PHI2X1(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X1),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X1_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1_number),
.read_add(VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1),
.start(PR_L5D3_L3L4_start),
.done(VMPROJ_L3L4_L5D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X1n5;
wire VMR_L5D3_VMS_L5D3PHI2X1n5_wr_en;
wire [5:0] VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1_number;
wire [10:0] VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1_read_add;
wire [18:0] VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1;
VMStubs #("Match") VMS_L5D3PHI2X1n5(
.data_in(VMR_L5D3_VMS_L5D3PHI2X1n5),
.enable(VMR_L5D3_VMS_L5D3PHI2X1n5_wr_en),
.number_out(VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1_number),
.read_add(VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1_read_add),
.data_out(VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X2;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2_read_add;
wire [13:0] VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2;
VMProjections  VMPROJ_L3L4_L5D3PHI2X2(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X2),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X2_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2_number),
.read_add(VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2),
.start(PR_L5D3_L3L4_start),
.done(VMPROJ_L3L4_L5D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X2n5;
wire VMR_L5D3_VMS_L5D3PHI2X2n5_wr_en;
wire [5:0] VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2_number;
wire [10:0] VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2_read_add;
wire [18:0] VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2;
VMStubs #("Match") VMS_L5D3PHI2X2n5(
.data_in(VMR_L5D3_VMS_L5D3PHI2X2n5),
.enable(VMR_L5D3_VMS_L5D3PHI2X2n5_wr_en),
.number_out(VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2_number),
.read_add(VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2_read_add),
.data_out(VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X1;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1_read_add;
wire [13:0] VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1;
VMProjections  VMPROJ_L3L4_L5D3PHI3X1(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X1),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X1_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1_number),
.read_add(VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1),
.start(PR_L5D3_L3L4_start),
.done(VMPROJ_L3L4_L5D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X1n5;
wire VMR_L5D3_VMS_L5D3PHI3X1n5_wr_en;
wire [5:0] VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1_number;
wire [10:0] VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1_read_add;
wire [18:0] VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1;
VMStubs #("Match") VMS_L5D3PHI3X1n5(
.data_in(VMR_L5D3_VMS_L5D3PHI3X1n5),
.enable(VMR_L5D3_VMS_L5D3PHI3X1n5_wr_en),
.number_out(VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1_number),
.read_add(VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1_read_add),
.data_out(VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X2;
wire PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2_number;
wire [8:0] VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2_read_add;
wire [13:0] VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2;
VMProjections  VMPROJ_L3L4_L5D3PHI3X2(
.data_in(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X2),
.enable(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X2_wr_en),
.number_out(VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2_number),
.read_add(VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2_read_add),
.data_out(VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2),
.start(PR_L5D3_L3L4_start),
.done(VMPROJ_L3L4_L5D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X2n5;
wire VMR_L5D3_VMS_L5D3PHI3X2n5_wr_en;
wire [5:0] VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2_number;
wire [10:0] VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2_read_add;
wire [18:0] VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2;
VMStubs #("Match") VMS_L5D3PHI3X2n5(
.data_in(VMR_L5D3_VMS_L5D3PHI3X2n5),
.enable(VMR_L5D3_VMS_L5D3PHI3X2n5_wr_en),
.number_out(VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2_number),
.read_add(VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2_read_add),
.data_out(VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X1;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1_read_add;
wire [13:0] VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1;
VMProjections  VMPROJ_L3L4_L5D4PHI1X1(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X1),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X1_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1_number),
.read_add(VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1),
.start(PR_L5D4_L3L4_start),
.done(VMPROJ_L3L4_L5D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X1n5;
wire VMR_L5D4_VMS_L5D4PHI1X1n5_wr_en;
wire [5:0] VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1_number;
wire [10:0] VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1_read_add;
wire [18:0] VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1;
VMStubs #("Match") VMS_L5D4PHI1X1n5(
.data_in(VMR_L5D4_VMS_L5D4PHI1X1n5),
.enable(VMR_L5D4_VMS_L5D4PHI1X1n5_wr_en),
.number_out(VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1_number),
.read_add(VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1_read_add),
.data_out(VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X2;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2_read_add;
wire [13:0] VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2;
VMProjections  VMPROJ_L3L4_L5D4PHI1X2(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X2),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X2_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2_number),
.read_add(VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2),
.start(PR_L5D4_L3L4_start),
.done(VMPROJ_L3L4_L5D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X2n3;
wire VMR_L5D4_VMS_L5D4PHI1X2n3_wr_en;
wire [5:0] VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2_number;
wire [10:0] VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2_read_add;
wire [18:0] VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2;
VMStubs #("Match") VMS_L5D4PHI1X2n3(
.data_in(VMR_L5D4_VMS_L5D4PHI1X2n3),
.enable(VMR_L5D4_VMS_L5D4PHI1X2n3_wr_en),
.number_out(VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2_number),
.read_add(VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2_read_add),
.data_out(VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X1;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1_read_add;
wire [13:0] VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1;
VMProjections  VMPROJ_L3L4_L5D4PHI2X1(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X1),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X1_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1_number),
.read_add(VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1),
.start(PR_L5D4_L3L4_start),
.done(VMPROJ_L3L4_L5D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X1n5;
wire VMR_L5D4_VMS_L5D4PHI2X1n5_wr_en;
wire [5:0] VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1_number;
wire [10:0] VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1_read_add;
wire [18:0] VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1;
VMStubs #("Match") VMS_L5D4PHI2X1n5(
.data_in(VMR_L5D4_VMS_L5D4PHI2X1n5),
.enable(VMR_L5D4_VMS_L5D4PHI2X1n5_wr_en),
.number_out(VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1_number),
.read_add(VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1_read_add),
.data_out(VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X2;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2_read_add;
wire [13:0] VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2;
VMProjections  VMPROJ_L3L4_L5D4PHI2X2(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X2),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X2_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2_number),
.read_add(VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2),
.start(PR_L5D4_L3L4_start),
.done(VMPROJ_L3L4_L5D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X2n3;
wire VMR_L5D4_VMS_L5D4PHI2X2n3_wr_en;
wire [5:0] VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2_number;
wire [10:0] VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2_read_add;
wire [18:0] VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2;
VMStubs #("Match") VMS_L5D4PHI2X2n3(
.data_in(VMR_L5D4_VMS_L5D4PHI2X2n3),
.enable(VMR_L5D4_VMS_L5D4PHI2X2n3_wr_en),
.number_out(VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2_number),
.read_add(VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2_read_add),
.data_out(VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X1;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1_read_add;
wire [13:0] VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1;
VMProjections  VMPROJ_L3L4_L5D4PHI3X1(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X1),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X1_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1_number),
.read_add(VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1),
.start(PR_L5D4_L3L4_start),
.done(VMPROJ_L3L4_L5D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X1n5;
wire VMR_L5D4_VMS_L5D4PHI3X1n5_wr_en;
wire [5:0] VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1_number;
wire [10:0] VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1_read_add;
wire [18:0] VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1;
VMStubs #("Match") VMS_L5D4PHI3X1n5(
.data_in(VMR_L5D4_VMS_L5D4PHI3X1n5),
.enable(VMR_L5D4_VMS_L5D4PHI3X1n5_wr_en),
.number_out(VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1_number),
.read_add(VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1_read_add),
.data_out(VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X2;
wire PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2_number;
wire [8:0] VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2_read_add;
wire [13:0] VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2;
VMProjections  VMPROJ_L3L4_L5D4PHI3X2(
.data_in(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X2),
.enable(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X2_wr_en),
.number_out(VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2_number),
.read_add(VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2_read_add),
.data_out(VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2),
.start(PR_L5D4_L3L4_start),
.done(VMPROJ_L3L4_L5D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X2n3;
wire VMR_L5D4_VMS_L5D4PHI3X2n3_wr_en;
wire [5:0] VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2_number;
wire [10:0] VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2_read_add;
wire [18:0] VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2;
VMStubs #("Match") VMS_L5D4PHI3X2n3(
.data_in(VMR_L5D4_VMS_L5D4PHI3X2n3),
.enable(VMR_L5D4_VMS_L5D4PHI3X2n3_wr_en),
.number_out(VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2_number),
.read_add(VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2_read_add),
.data_out(VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X1;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1_read_add;
wire [13:0] VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1;
VMProjections  VMPROJ_L3L4_L6D3PHI1X1(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X1),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X1_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1_number),
.read_add(VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1),
.start(PR_L6D3_L3L4_start),
.done(VMPROJ_L3L4_L6D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI1X1n2;
wire VMR_L6D3_VMS_L6D3PHI1X1n2_wr_en;
wire [5:0] VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1_number;
wire [10:0] VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1_read_add;
wire [18:0] VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1;
VMStubs #("Match") VMS_L6D3PHI1X1n2(
.data_in(VMR_L6D3_VMS_L6D3PHI1X1n2),
.enable(VMR_L6D3_VMS_L6D3PHI1X1n2_wr_en),
.number_out(VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1_number),
.read_add(VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1_read_add),
.data_out(VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X2;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2_read_add;
wire [13:0] VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2;
VMProjections  VMPROJ_L3L4_L6D3PHI1X2(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X2),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X2_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2_number),
.read_add(VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2),
.start(PR_L6D3_L3L4_start),
.done(VMPROJ_L3L4_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI1X2n3;
wire VMR_L6D3_VMS_L6D3PHI1X2n3_wr_en;
wire [5:0] VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2_number;
wire [10:0] VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2_read_add;
wire [18:0] VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2;
VMStubs #("Match") VMS_L6D3PHI1X2n3(
.data_in(VMR_L6D3_VMS_L6D3PHI1X2n3),
.enable(VMR_L6D3_VMS_L6D3PHI1X2n3_wr_en),
.number_out(VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2_number),
.read_add(VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2_read_add),
.data_out(VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X1;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1_read_add;
wire [13:0] VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1;
VMProjections  VMPROJ_L3L4_L6D3PHI2X1(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X1),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X1_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1_number),
.read_add(VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1),
.start(PR_L6D3_L3L4_start),
.done(VMPROJ_L3L4_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X1n3;
wire VMR_L6D3_VMS_L6D3PHI2X1n3_wr_en;
wire [5:0] VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1_number;
wire [10:0] VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1_read_add;
wire [18:0] VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1;
VMStubs #("Match") VMS_L6D3PHI2X1n3(
.data_in(VMR_L6D3_VMS_L6D3PHI2X1n3),
.enable(VMR_L6D3_VMS_L6D3PHI2X1n3_wr_en),
.number_out(VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1_number),
.read_add(VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1_read_add),
.data_out(VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X2;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2_read_add;
wire [13:0] VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2;
VMProjections  VMPROJ_L3L4_L6D3PHI2X2(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X2),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X2_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2_number),
.read_add(VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2),
.start(PR_L6D3_L3L4_start),
.done(VMPROJ_L3L4_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X2n5;
wire VMR_L6D3_VMS_L6D3PHI2X2n5_wr_en;
wire [5:0] VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2_number;
wire [10:0] VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2_read_add;
wire [18:0] VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2;
VMStubs #("Match") VMS_L6D3PHI2X2n5(
.data_in(VMR_L6D3_VMS_L6D3PHI2X2n5),
.enable(VMR_L6D3_VMS_L6D3PHI2X2n5_wr_en),
.number_out(VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2_number),
.read_add(VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2_read_add),
.data_out(VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X1;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1_read_add;
wire [13:0] VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1;
VMProjections  VMPROJ_L3L4_L6D3PHI3X1(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X1),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X1_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1_number),
.read_add(VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1),
.start(PR_L6D3_L3L4_start),
.done(VMPROJ_L3L4_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X1n3;
wire VMR_L6D3_VMS_L6D3PHI3X1n3_wr_en;
wire [5:0] VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1_number;
wire [10:0] VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1_read_add;
wire [18:0] VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1;
VMStubs #("Match") VMS_L6D3PHI3X1n3(
.data_in(VMR_L6D3_VMS_L6D3PHI3X1n3),
.enable(VMR_L6D3_VMS_L6D3PHI3X1n3_wr_en),
.number_out(VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1_number),
.read_add(VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1_read_add),
.data_out(VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X2;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2_read_add;
wire [13:0] VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2;
VMProjections  VMPROJ_L3L4_L6D3PHI3X2(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X2),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X2_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2_number),
.read_add(VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2),
.start(PR_L6D3_L3L4_start),
.done(VMPROJ_L3L4_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X2n5;
wire VMR_L6D3_VMS_L6D3PHI3X2n5_wr_en;
wire [5:0] VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2_number;
wire [10:0] VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2_read_add;
wire [18:0] VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2;
VMStubs #("Match") VMS_L6D3PHI3X2n5(
.data_in(VMR_L6D3_VMS_L6D3PHI3X2n5),
.enable(VMR_L6D3_VMS_L6D3PHI3X2n5_wr_en),
.number_out(VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2_number),
.read_add(VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2_read_add),
.data_out(VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X1;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1_read_add;
wire [13:0] VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1;
VMProjections  VMPROJ_L3L4_L6D3PHI4X1(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X1),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X1_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1_number),
.read_add(VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1),
.start(PR_L6D3_L3L4_start),
.done(VMPROJ_L3L4_L6D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI4X1n2;
wire VMR_L6D3_VMS_L6D3PHI4X1n2_wr_en;
wire [5:0] VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1_number;
wire [10:0] VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1_read_add;
wire [18:0] VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1;
VMStubs #("Match") VMS_L6D3PHI4X1n2(
.data_in(VMR_L6D3_VMS_L6D3PHI4X1n2),
.enable(VMR_L6D3_VMS_L6D3PHI4X1n2_wr_en),
.number_out(VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1_number),
.read_add(VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1_read_add),
.data_out(VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X2;
wire PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2_number;
wire [8:0] VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2_read_add;
wire [13:0] VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2;
VMProjections  VMPROJ_L3L4_L6D3PHI4X2(
.data_in(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X2),
.enable(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X2_wr_en),
.number_out(VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2_number),
.read_add(VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2_read_add),
.data_out(VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2),
.start(PR_L6D3_L3L4_start),
.done(VMPROJ_L3L4_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI4X2n3;
wire VMR_L6D3_VMS_L6D3PHI4X2n3_wr_en;
wire [5:0] VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2_number;
wire [10:0] VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2_read_add;
wire [18:0] VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2;
VMStubs #("Match") VMS_L6D3PHI4X2n3(
.data_in(VMR_L6D3_VMS_L6D3PHI4X2n3),
.enable(VMR_L6D3_VMS_L6D3PHI4X2n3_wr_en),
.number_out(VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2_number),
.read_add(VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2_read_add),
.data_out(VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI4X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X1;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1_read_add;
wire [13:0] VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1;
VMProjections  VMPROJ_L3L4_L6D4PHI1X1(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X1),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X1_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1_number),
.read_add(VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1),
.start(PR_L6D4_L3L4_start),
.done(VMPROJ_L3L4_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI1X1n3;
wire VMR_L6D4_VMS_L6D4PHI1X1n3_wr_en;
wire [5:0] VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1_number;
wire [10:0] VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1_read_add;
wire [18:0] VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1;
VMStubs #("Match") VMS_L6D4PHI1X1n3(
.data_in(VMR_L6D4_VMS_L6D4PHI1X1n3),
.enable(VMR_L6D4_VMS_L6D4PHI1X1n3_wr_en),
.number_out(VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1_number),
.read_add(VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1_read_add),
.data_out(VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X2;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2_read_add;
wire [13:0] VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2;
VMProjections  VMPROJ_L3L4_L6D4PHI1X2(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X2),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X2_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2_number),
.read_add(VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2),
.start(PR_L6D4_L3L4_start),
.done(VMPROJ_L3L4_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI1X2n3;
wire VMR_L6D4_VMS_L6D4PHI1X2n3_wr_en;
wire [5:0] VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2_number;
wire [10:0] VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2_read_add;
wire [18:0] VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2;
VMStubs #("Match") VMS_L6D4PHI1X2n3(
.data_in(VMR_L6D4_VMS_L6D4PHI1X2n3),
.enable(VMR_L6D4_VMS_L6D4PHI1X2n3_wr_en),
.number_out(VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2_number),
.read_add(VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2_read_add),
.data_out(VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X1;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1_read_add;
wire [13:0] VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1;
VMProjections  VMPROJ_L3L4_L6D4PHI2X1(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X1),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X1_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1_number),
.read_add(VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1),
.start(PR_L6D4_L3L4_start),
.done(VMPROJ_L3L4_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X1n5;
wire VMR_L6D4_VMS_L6D4PHI2X1n5_wr_en;
wire [5:0] VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1_number;
wire [10:0] VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1_read_add;
wire [18:0] VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1;
VMStubs #("Match") VMS_L6D4PHI2X1n5(
.data_in(VMR_L6D4_VMS_L6D4PHI2X1n5),
.enable(VMR_L6D4_VMS_L6D4PHI2X1n5_wr_en),
.number_out(VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1_number),
.read_add(VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1_read_add),
.data_out(VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X2;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2_read_add;
wire [13:0] VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2;
VMProjections  VMPROJ_L3L4_L6D4PHI2X2(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X2),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X2_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2_number),
.read_add(VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2),
.start(PR_L6D4_L3L4_start),
.done(VMPROJ_L3L4_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X2n5;
wire VMR_L6D4_VMS_L6D4PHI2X2n5_wr_en;
wire [5:0] VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2_number;
wire [10:0] VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2_read_add;
wire [18:0] VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2;
VMStubs #("Match") VMS_L6D4PHI2X2n5(
.data_in(VMR_L6D4_VMS_L6D4PHI2X2n5),
.enable(VMR_L6D4_VMS_L6D4PHI2X2n5_wr_en),
.number_out(VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2_number),
.read_add(VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2_read_add),
.data_out(VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X1;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1_read_add;
wire [13:0] VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1;
VMProjections  VMPROJ_L3L4_L6D4PHI3X1(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X1),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X1_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1_number),
.read_add(VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1),
.start(PR_L6D4_L3L4_start),
.done(VMPROJ_L3L4_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X1n5;
wire VMR_L6D4_VMS_L6D4PHI3X1n5_wr_en;
wire [5:0] VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1_number;
wire [10:0] VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1_read_add;
wire [18:0] VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1;
VMStubs #("Match") VMS_L6D4PHI3X1n5(
.data_in(VMR_L6D4_VMS_L6D4PHI3X1n5),
.enable(VMR_L6D4_VMS_L6D4PHI3X1n5_wr_en),
.number_out(VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1_number),
.read_add(VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1_read_add),
.data_out(VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X2;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2_read_add;
wire [13:0] VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2;
VMProjections  VMPROJ_L3L4_L6D4PHI3X2(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X2),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X2_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2_number),
.read_add(VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2),
.start(PR_L6D4_L3L4_start),
.done(VMPROJ_L3L4_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X2n5;
wire VMR_L6D4_VMS_L6D4PHI3X2n5_wr_en;
wire [5:0] VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2_number;
wire [10:0] VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2_read_add;
wire [18:0] VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2;
VMStubs #("Match") VMS_L6D4PHI3X2n5(
.data_in(VMR_L6D4_VMS_L6D4PHI3X2n5),
.enable(VMR_L6D4_VMS_L6D4PHI3X2n5_wr_en),
.number_out(VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2_number),
.read_add(VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2_read_add),
.data_out(VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X1;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X1_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1_read_add;
wire [13:0] VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1;
VMProjections  VMPROJ_L3L4_L6D4PHI4X1(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X1),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X1_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1_number),
.read_add(VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1),
.start(PR_L6D4_L3L4_start),
.done(VMPROJ_L3L4_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI4X1n3;
wire VMR_L6D4_VMS_L6D4PHI4X1n3_wr_en;
wire [5:0] VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1_number;
wire [10:0] VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1_read_add;
wire [18:0] VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1;
VMStubs #("Match") VMS_L6D4PHI4X1n3(
.data_in(VMR_L6D4_VMS_L6D4PHI4X1n3),
.enable(VMR_L6D4_VMS_L6D4PHI4X1n3_wr_en),
.number_out(VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1_number),
.read_add(VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1_read_add),
.data_out(VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI4X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X2;
wire PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X2_wr_en;
wire [5:0] VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2_number;
wire [8:0] VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2_read_add;
wire [13:0] VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2;
VMProjections  VMPROJ_L3L4_L6D4PHI4X2(
.data_in(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X2),
.enable(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X2_wr_en),
.number_out(VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2_number),
.read_add(VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2_read_add),
.data_out(VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2),
.start(PR_L6D4_L3L4_start),
.done(VMPROJ_L3L4_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI4X2n3;
wire VMR_L6D4_VMS_L6D4PHI4X2n3_wr_en;
wire [5:0] VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2_number;
wire [10:0] VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2_read_add;
wire [18:0] VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2;
VMStubs #("Match") VMS_L6D4PHI4X2n3(
.data_in(VMR_L6D4_VMS_L6D4PHI4X2n3),
.enable(VMR_L6D4_VMS_L6D4PHI4X2n3_wr_en),
.number_out(VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2_number),
.read_add(VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2_read_add),
.data_out(VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI4X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X1;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1_read_add;
wire [13:0] VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1;
VMProjections  VMPROJ_L1L2_L3D3PHI1X1(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X1),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X1_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1_number),
.read_add(VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1),
.start(PR_L3D3_L1L2_start),
.done(VMPROJ_L1L2_L3D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X1n5;
wire VMR_L3D3_VMS_L3D3PHI1X1n5_wr_en;
wire [5:0] VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1_number;
wire [10:0] VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1_read_add;
wire [18:0] VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1;
VMStubs #("Match") VMS_L3D3PHI1X1n5(
.data_in(VMR_L3D3_VMS_L3D3PHI1X1n5),
.enable(VMR_L3D3_VMS_L3D3PHI1X1n5_wr_en),
.number_out(VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1_number),
.read_add(VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1_read_add),
.data_out(VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X2;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2_read_add;
wire [13:0] VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2;
VMProjections  VMPROJ_L1L2_L3D3PHI1X2(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X2),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X2_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2_number),
.read_add(VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2),
.start(PR_L3D3_L1L2_start),
.done(VMPROJ_L1L2_L3D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X2n5;
wire VMR_L3D3_VMS_L3D3PHI1X2n5_wr_en;
wire [5:0] VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2_number;
wire [10:0] VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2_read_add;
wire [18:0] VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2;
VMStubs #("Match") VMS_L3D3PHI1X2n5(
.data_in(VMR_L3D3_VMS_L3D3PHI1X2n5),
.enable(VMR_L3D3_VMS_L3D3PHI1X2n5_wr_en),
.number_out(VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2_number),
.read_add(VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2_read_add),
.data_out(VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X1;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1_read_add;
wire [13:0] VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1;
VMProjections  VMPROJ_L1L2_L3D3PHI2X1(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X1),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X1_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1_number),
.read_add(VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1),
.start(PR_L3D3_L1L2_start),
.done(VMPROJ_L1L2_L3D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X1n5;
wire VMR_L3D3_VMS_L3D3PHI2X1n5_wr_en;
wire [5:0] VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1_number;
wire [10:0] VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1_read_add;
wire [18:0] VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1;
VMStubs #("Match") VMS_L3D3PHI2X1n5(
.data_in(VMR_L3D3_VMS_L3D3PHI2X1n5),
.enable(VMR_L3D3_VMS_L3D3PHI2X1n5_wr_en),
.number_out(VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1_number),
.read_add(VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1_read_add),
.data_out(VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X2;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2_read_add;
wire [13:0] VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2;
VMProjections  VMPROJ_L1L2_L3D3PHI2X2(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X2),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X2_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2_number),
.read_add(VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2),
.start(PR_L3D3_L1L2_start),
.done(VMPROJ_L1L2_L3D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X2n5;
wire VMR_L3D3_VMS_L3D3PHI2X2n5_wr_en;
wire [5:0] VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2_number;
wire [10:0] VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2_read_add;
wire [18:0] VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2;
VMStubs #("Match") VMS_L3D3PHI2X2n5(
.data_in(VMR_L3D3_VMS_L3D3PHI2X2n5),
.enable(VMR_L3D3_VMS_L3D3PHI2X2n5_wr_en),
.number_out(VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2_number),
.read_add(VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2_read_add),
.data_out(VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X1;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1_read_add;
wire [13:0] VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1;
VMProjections  VMPROJ_L1L2_L3D3PHI3X1(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X1),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X1_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1_number),
.read_add(VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1),
.start(PR_L3D3_L1L2_start),
.done(VMPROJ_L1L2_L3D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X1n5;
wire VMR_L3D3_VMS_L3D3PHI3X1n5_wr_en;
wire [5:0] VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1_number;
wire [10:0] VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1_read_add;
wire [18:0] VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1;
VMStubs #("Match") VMS_L3D3PHI3X1n5(
.data_in(VMR_L3D3_VMS_L3D3PHI3X1n5),
.enable(VMR_L3D3_VMS_L3D3PHI3X1n5_wr_en),
.number_out(VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1_number),
.read_add(VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1_read_add),
.data_out(VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X2;
wire PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2_number;
wire [8:0] VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2_read_add;
wire [13:0] VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2;
VMProjections  VMPROJ_L1L2_L3D3PHI3X2(
.data_in(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X2),
.enable(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X2_wr_en),
.number_out(VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2_number),
.read_add(VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2_read_add),
.data_out(VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2),
.start(PR_L3D3_L1L2_start),
.done(VMPROJ_L1L2_L3D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X2n5;
wire VMR_L3D3_VMS_L3D3PHI3X2n5_wr_en;
wire [5:0] VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2_number;
wire [10:0] VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2_read_add;
wire [18:0] VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2;
VMStubs #("Match") VMS_L3D3PHI3X2n5(
.data_in(VMR_L3D3_VMS_L3D3PHI3X2n5),
.enable(VMR_L3D3_VMS_L3D3PHI3X2n5_wr_en),
.number_out(VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2_number),
.read_add(VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2_read_add),
.data_out(VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X1;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1_read_add;
wire [13:0] VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1;
VMProjections  VMPROJ_L1L2_L3D4PHI1X1(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X1),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X1_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1_number),
.read_add(VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1),
.start(PR_L3D4_L1L2_start),
.done(VMPROJ_L1L2_L3D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X1n5;
wire VMR_L3D4_VMS_L3D4PHI1X1n5_wr_en;
wire [5:0] VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1_number;
wire [10:0] VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1_read_add;
wire [18:0] VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1;
VMStubs #("Match") VMS_L3D4PHI1X1n5(
.data_in(VMR_L3D4_VMS_L3D4PHI1X1n5),
.enable(VMR_L3D4_VMS_L3D4PHI1X1n5_wr_en),
.number_out(VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1_number),
.read_add(VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1_read_add),
.data_out(VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X2;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2_read_add;
wire [13:0] VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2;
VMProjections  VMPROJ_L1L2_L3D4PHI1X2(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X2),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X2_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2_number),
.read_add(VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2),
.start(PR_L3D4_L1L2_start),
.done(VMPROJ_L1L2_L3D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X2n3;
wire VMR_L3D4_VMS_L3D4PHI1X2n3_wr_en;
wire [5:0] VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2_number;
wire [10:0] VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2_read_add;
wire [18:0] VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2;
VMStubs #("Match") VMS_L3D4PHI1X2n3(
.data_in(VMR_L3D4_VMS_L3D4PHI1X2n3),
.enable(VMR_L3D4_VMS_L3D4PHI1X2n3_wr_en),
.number_out(VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2_number),
.read_add(VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2_read_add),
.data_out(VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X1;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1_read_add;
wire [13:0] VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1;
VMProjections  VMPROJ_L1L2_L3D4PHI2X1(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X1),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X1_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1_number),
.read_add(VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1),
.start(PR_L3D4_L1L2_start),
.done(VMPROJ_L1L2_L3D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X1n5;
wire VMR_L3D4_VMS_L3D4PHI2X1n5_wr_en;
wire [5:0] VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1_number;
wire [10:0] VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1_read_add;
wire [18:0] VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1;
VMStubs #("Match") VMS_L3D4PHI2X1n5(
.data_in(VMR_L3D4_VMS_L3D4PHI2X1n5),
.enable(VMR_L3D4_VMS_L3D4PHI2X1n5_wr_en),
.number_out(VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1_number),
.read_add(VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1_read_add),
.data_out(VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X2;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2_read_add;
wire [13:0] VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2;
VMProjections  VMPROJ_L1L2_L3D4PHI2X2(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X2),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X2_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2_number),
.read_add(VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2),
.start(PR_L3D4_L1L2_start),
.done(VMPROJ_L1L2_L3D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X2n3;
wire VMR_L3D4_VMS_L3D4PHI2X2n3_wr_en;
wire [5:0] VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2_number;
wire [10:0] VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2_read_add;
wire [18:0] VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2;
VMStubs #("Match") VMS_L3D4PHI2X2n3(
.data_in(VMR_L3D4_VMS_L3D4PHI2X2n3),
.enable(VMR_L3D4_VMS_L3D4PHI2X2n3_wr_en),
.number_out(VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2_number),
.read_add(VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2_read_add),
.data_out(VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X1;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1_read_add;
wire [13:0] VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1;
VMProjections  VMPROJ_L1L2_L3D4PHI3X1(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X1),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X1_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1_number),
.read_add(VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1),
.start(PR_L3D4_L1L2_start),
.done(VMPROJ_L1L2_L3D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X1n5;
wire VMR_L3D4_VMS_L3D4PHI3X1n5_wr_en;
wire [5:0] VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1_number;
wire [10:0] VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1_read_add;
wire [18:0] VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1;
VMStubs #("Match") VMS_L3D4PHI3X1n5(
.data_in(VMR_L3D4_VMS_L3D4PHI3X1n5),
.enable(VMR_L3D4_VMS_L3D4PHI3X1n5_wr_en),
.number_out(VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1_number),
.read_add(VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1_read_add),
.data_out(VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X2;
wire PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2_number;
wire [8:0] VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2_read_add;
wire [13:0] VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2;
VMProjections  VMPROJ_L1L2_L3D4PHI3X2(
.data_in(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X2),
.enable(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X2_wr_en),
.number_out(VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2_number),
.read_add(VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2_read_add),
.data_out(VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2),
.start(PR_L3D4_L1L2_start),
.done(VMPROJ_L1L2_L3D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X2n3;
wire VMR_L3D4_VMS_L3D4PHI3X2n3_wr_en;
wire [5:0] VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2_number;
wire [10:0] VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2_read_add;
wire [18:0] VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2;
VMStubs #("Match") VMS_L3D4PHI3X2n3(
.data_in(VMR_L3D4_VMS_L3D4PHI3X2n3),
.enable(VMR_L3D4_VMS_L3D4PHI3X2n3_wr_en),
.number_out(VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2_number),
.read_add(VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2_read_add),
.data_out(VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X1;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1_read_add;
wire [13:0] VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1;
VMProjections  VMPROJ_L1L2_L4D3PHI1X1(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X1),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X1_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1_number),
.read_add(VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1),
.start(PR_L4D3_L1L2_start),
.done(VMPROJ_L1L2_L4D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI1X1n2;
wire VMR_L4D3_VMS_L4D3PHI1X1n2_wr_en;
wire [5:0] VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1_number;
wire [10:0] VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1_read_add;
wire [18:0] VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1;
VMStubs #("Match") VMS_L4D3PHI1X1n2(
.data_in(VMR_L4D3_VMS_L4D3PHI1X1n2),
.enable(VMR_L4D3_VMS_L4D3PHI1X1n2_wr_en),
.number_out(VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1_number),
.read_add(VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1_read_add),
.data_out(VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI1X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X2;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2_read_add;
wire [13:0] VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2;
VMProjections  VMPROJ_L1L2_L4D3PHI1X2(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X2),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X2_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2_number),
.read_add(VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2),
.start(PR_L4D3_L1L2_start),
.done(VMPROJ_L1L2_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI1X2n3;
wire VMR_L4D3_VMS_L4D3PHI1X2n3_wr_en;
wire [5:0] VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2_number;
wire [10:0] VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2_read_add;
wire [18:0] VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2;
VMStubs #("Match") VMS_L4D3PHI1X2n3(
.data_in(VMR_L4D3_VMS_L4D3PHI1X2n3),
.enable(VMR_L4D3_VMS_L4D3PHI1X2n3_wr_en),
.number_out(VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2_number),
.read_add(VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2_read_add),
.data_out(VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X1;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1_read_add;
wire [13:0] VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1;
VMProjections  VMPROJ_L1L2_L4D3PHI2X1(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X1),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X1_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1_number),
.read_add(VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1),
.start(PR_L4D3_L1L2_start),
.done(VMPROJ_L1L2_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X1n3;
wire VMR_L4D3_VMS_L4D3PHI2X1n3_wr_en;
wire [5:0] VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1_number;
wire [10:0] VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1_read_add;
wire [18:0] VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1;
VMStubs #("Match") VMS_L4D3PHI2X1n3(
.data_in(VMR_L4D3_VMS_L4D3PHI2X1n3),
.enable(VMR_L4D3_VMS_L4D3PHI2X1n3_wr_en),
.number_out(VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1_number),
.read_add(VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1_read_add),
.data_out(VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X2;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2_read_add;
wire [13:0] VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2;
VMProjections  VMPROJ_L1L2_L4D3PHI2X2(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X2),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X2_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2_number),
.read_add(VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2),
.start(PR_L4D3_L1L2_start),
.done(VMPROJ_L1L2_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X2n5;
wire VMR_L4D3_VMS_L4D3PHI2X2n5_wr_en;
wire [5:0] VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2_number;
wire [10:0] VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2_read_add;
wire [18:0] VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2;
VMStubs #("Match") VMS_L4D3PHI2X2n5(
.data_in(VMR_L4D3_VMS_L4D3PHI2X2n5),
.enable(VMR_L4D3_VMS_L4D3PHI2X2n5_wr_en),
.number_out(VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2_number),
.read_add(VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2_read_add),
.data_out(VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X1;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1_read_add;
wire [13:0] VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1;
VMProjections  VMPROJ_L1L2_L4D3PHI3X1(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X1),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X1_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1_number),
.read_add(VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1),
.start(PR_L4D3_L1L2_start),
.done(VMPROJ_L1L2_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X1n3;
wire VMR_L4D3_VMS_L4D3PHI3X1n3_wr_en;
wire [5:0] VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1_number;
wire [10:0] VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1_read_add;
wire [18:0] VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1;
VMStubs #("Match") VMS_L4D3PHI3X1n3(
.data_in(VMR_L4D3_VMS_L4D3PHI3X1n3),
.enable(VMR_L4D3_VMS_L4D3PHI3X1n3_wr_en),
.number_out(VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1_number),
.read_add(VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1_read_add),
.data_out(VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X2;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2_read_add;
wire [13:0] VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2;
VMProjections  VMPROJ_L1L2_L4D3PHI3X2(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X2),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X2_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2_number),
.read_add(VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2),
.start(PR_L4D3_L1L2_start),
.done(VMPROJ_L1L2_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X2n5;
wire VMR_L4D3_VMS_L4D3PHI3X2n5_wr_en;
wire [5:0] VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2_number;
wire [10:0] VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2_read_add;
wire [18:0] VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2;
VMStubs #("Match") VMS_L4D3PHI3X2n5(
.data_in(VMR_L4D3_VMS_L4D3PHI3X2n5),
.enable(VMR_L4D3_VMS_L4D3PHI3X2n5_wr_en),
.number_out(VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2_number),
.read_add(VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2_read_add),
.data_out(VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X1;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1_read_add;
wire [13:0] VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1;
VMProjections  VMPROJ_L1L2_L4D3PHI4X1(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X1),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X1_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1_number),
.read_add(VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1),
.start(PR_L4D3_L1L2_start),
.done(VMPROJ_L1L2_L4D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI4X1n2;
wire VMR_L4D3_VMS_L4D3PHI4X1n2_wr_en;
wire [5:0] VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1_number;
wire [10:0] VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1_read_add;
wire [18:0] VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1;
VMStubs #("Match") VMS_L4D3PHI4X1n2(
.data_in(VMR_L4D3_VMS_L4D3PHI4X1n2),
.enable(VMR_L4D3_VMS_L4D3PHI4X1n2_wr_en),
.number_out(VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1_number),
.read_add(VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1_read_add),
.data_out(VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI4X1n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X2;
wire PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2_number;
wire [8:0] VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2_read_add;
wire [13:0] VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2;
VMProjections  VMPROJ_L1L2_L4D3PHI4X2(
.data_in(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X2),
.enable(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X2_wr_en),
.number_out(VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2_number),
.read_add(VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2_read_add),
.data_out(VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2),
.start(PR_L4D3_L1L2_start),
.done(VMPROJ_L1L2_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI4X2n3;
wire VMR_L4D3_VMS_L4D3PHI4X2n3_wr_en;
wire [5:0] VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2_number;
wire [10:0] VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2_read_add;
wire [18:0] VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2;
VMStubs #("Match") VMS_L4D3PHI4X2n3(
.data_in(VMR_L4D3_VMS_L4D3PHI4X2n3),
.enable(VMR_L4D3_VMS_L4D3PHI4X2n3_wr_en),
.number_out(VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2_number),
.read_add(VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2_read_add),
.data_out(VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI4X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X1;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1_read_add;
wire [13:0] VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1;
VMProjections  VMPROJ_L1L2_L4D4PHI1X1(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X1),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X1_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1_number),
.read_add(VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1),
.start(PR_L4D4_L1L2_start),
.done(VMPROJ_L1L2_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI1X1n3;
wire VMR_L4D4_VMS_L4D4PHI1X1n3_wr_en;
wire [5:0] VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1_number;
wire [10:0] VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1_read_add;
wire [18:0] VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1;
VMStubs #("Match") VMS_L4D4PHI1X1n3(
.data_in(VMR_L4D4_VMS_L4D4PHI1X1n3),
.enable(VMR_L4D4_VMS_L4D4PHI1X1n3_wr_en),
.number_out(VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1_number),
.read_add(VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1_read_add),
.data_out(VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X2;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2_read_add;
wire [13:0] VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2;
VMProjections  VMPROJ_L1L2_L4D4PHI1X2(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X2),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X2_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2_number),
.read_add(VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2),
.start(PR_L4D4_L1L2_start),
.done(VMPROJ_L1L2_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI1X2n3;
wire VMR_L4D4_VMS_L4D4PHI1X2n3_wr_en;
wire [5:0] VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2_number;
wire [10:0] VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2_read_add;
wire [18:0] VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2;
VMStubs #("Match") VMS_L4D4PHI1X2n3(
.data_in(VMR_L4D4_VMS_L4D4PHI1X2n3),
.enable(VMR_L4D4_VMS_L4D4PHI1X2n3_wr_en),
.number_out(VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2_number),
.read_add(VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2_read_add),
.data_out(VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI1X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X1;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1_read_add;
wire [13:0] VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1;
VMProjections  VMPROJ_L1L2_L4D4PHI2X1(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X1),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X1_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1_number),
.read_add(VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1),
.start(PR_L4D4_L1L2_start),
.done(VMPROJ_L1L2_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X1n5;
wire VMR_L4D4_VMS_L4D4PHI2X1n5_wr_en;
wire [5:0] VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1_number;
wire [10:0] VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1_read_add;
wire [18:0] VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1;
VMStubs #("Match") VMS_L4D4PHI2X1n5(
.data_in(VMR_L4D4_VMS_L4D4PHI2X1n5),
.enable(VMR_L4D4_VMS_L4D4PHI2X1n5_wr_en),
.number_out(VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1_number),
.read_add(VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1_read_add),
.data_out(VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X2;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2_read_add;
wire [13:0] VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2;
VMProjections  VMPROJ_L1L2_L4D4PHI2X2(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X2),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X2_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2_number),
.read_add(VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2),
.start(PR_L4D4_L1L2_start),
.done(VMPROJ_L1L2_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X2n5;
wire VMR_L4D4_VMS_L4D4PHI2X2n5_wr_en;
wire [5:0] VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2_number;
wire [10:0] VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2_read_add;
wire [18:0] VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2;
VMStubs #("Match") VMS_L4D4PHI2X2n5(
.data_in(VMR_L4D4_VMS_L4D4PHI2X2n5),
.enable(VMR_L4D4_VMS_L4D4PHI2X2n5_wr_en),
.number_out(VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2_number),
.read_add(VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2_read_add),
.data_out(VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X1;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1_read_add;
wire [13:0] VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1;
VMProjections  VMPROJ_L1L2_L4D4PHI3X1(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X1),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X1_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1_number),
.read_add(VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1),
.start(PR_L4D4_L1L2_start),
.done(VMPROJ_L1L2_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X1n5;
wire VMR_L4D4_VMS_L4D4PHI3X1n5_wr_en;
wire [5:0] VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1_number;
wire [10:0] VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1_read_add;
wire [18:0] VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1;
VMStubs #("Match") VMS_L4D4PHI3X1n5(
.data_in(VMR_L4D4_VMS_L4D4PHI3X1n5),
.enable(VMR_L4D4_VMS_L4D4PHI3X1n5_wr_en),
.number_out(VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1_number),
.read_add(VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1_read_add),
.data_out(VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X1n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X2;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2_read_add;
wire [13:0] VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2;
VMProjections  VMPROJ_L1L2_L4D4PHI3X2(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X2),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X2_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2_number),
.read_add(VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2),
.start(PR_L4D4_L1L2_start),
.done(VMPROJ_L1L2_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X2n5;
wire VMR_L4D4_VMS_L4D4PHI3X2n5_wr_en;
wire [5:0] VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2_number;
wire [10:0] VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2_read_add;
wire [18:0] VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2;
VMStubs #("Match") VMS_L4D4PHI3X2n5(
.data_in(VMR_L4D4_VMS_L4D4PHI3X2n5),
.enable(VMR_L4D4_VMS_L4D4PHI3X2n5_wr_en),
.number_out(VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2_number),
.read_add(VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2_read_add),
.data_out(VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X2n5_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X1;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X1_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1_read_add;
wire [13:0] VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1;
VMProjections  VMPROJ_L1L2_L4D4PHI4X1(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X1),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X1_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1_number),
.read_add(VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1),
.start(PR_L4D4_L1L2_start),
.done(VMPROJ_L1L2_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI4X1n3;
wire VMR_L4D4_VMS_L4D4PHI4X1n3_wr_en;
wire [5:0] VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1_number;
wire [10:0] VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1_read_add;
wire [18:0] VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1;
VMStubs #("Match") VMS_L4D4PHI4X1n3(
.data_in(VMR_L4D4_VMS_L4D4PHI4X1n3),
.enable(VMR_L4D4_VMS_L4D4PHI4X1n3_wr_en),
.number_out(VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1_number),
.read_add(VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1_read_add),
.data_out(VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI4X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X2;
wire PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X2_wr_en;
wire [5:0] VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2_number;
wire [8:0] VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2_read_add;
wire [13:0] VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2;
VMProjections  VMPROJ_L1L2_L4D4PHI4X2(
.data_in(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X2),
.enable(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X2_wr_en),
.number_out(VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2_number),
.read_add(VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2_read_add),
.data_out(VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2),
.start(PR_L4D4_L1L2_start),
.done(VMPROJ_L1L2_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI4X2n3;
wire VMR_L4D4_VMS_L4D4PHI4X2n3_wr_en;
wire [5:0] VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2_number;
wire [10:0] VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2_read_add;
wire [18:0] VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2;
VMStubs #("Match") VMS_L4D4PHI4X2n3(
.data_in(VMR_L4D4_VMS_L4D4PHI4X2n3),
.enable(VMR_L4D4_VMS_L4D4PHI4X2n3_wr_en),
.number_out(VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2_number),
.read_add(VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2_read_add),
.data_out(VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI4X2n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X1;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1_read_add;
wire [13:0] VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1;
VMProjections  VMPROJ_L1L2_L5D3PHI1X1(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X1),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X1_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1_number),
.read_add(VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1),
.start(PR_L5D3_L1L2_start),
.done(VMPROJ_L1L2_L5D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X1n6;
wire VMR_L5D3_VMS_L5D3PHI1X1n6_wr_en;
wire [5:0] VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1_number;
wire [10:0] VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1_read_add;
wire [18:0] VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1;
VMStubs #("Match") VMS_L5D3PHI1X1n6(
.data_in(VMR_L5D3_VMS_L5D3PHI1X1n6),
.enable(VMR_L5D3_VMS_L5D3PHI1X1n6_wr_en),
.number_out(VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1_number),
.read_add(VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1_read_add),
.data_out(VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X2;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2_read_add;
wire [13:0] VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2;
VMProjections  VMPROJ_L1L2_L5D3PHI1X2(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X2),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X2_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2_number),
.read_add(VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2),
.start(PR_L5D3_L1L2_start),
.done(VMPROJ_L1L2_L5D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI1X2n6;
wire VMR_L5D3_VMS_L5D3PHI1X2n6_wr_en;
wire [5:0] VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2_number;
wire [10:0] VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2_read_add;
wire [18:0] VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2;
VMStubs #("Match") VMS_L5D3PHI1X2n6(
.data_in(VMR_L5D3_VMS_L5D3PHI1X2n6),
.enable(VMR_L5D3_VMS_L5D3PHI1X2n6_wr_en),
.number_out(VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2_number),
.read_add(VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2_read_add),
.data_out(VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI1X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X1;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1_read_add;
wire [13:0] VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1;
VMProjections  VMPROJ_L1L2_L5D3PHI2X1(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X1),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X1_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1_number),
.read_add(VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1),
.start(PR_L5D3_L1L2_start),
.done(VMPROJ_L1L2_L5D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X1n6;
wire VMR_L5D3_VMS_L5D3PHI2X1n6_wr_en;
wire [5:0] VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1_number;
wire [10:0] VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1_read_add;
wire [18:0] VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1;
VMStubs #("Match") VMS_L5D3PHI2X1n6(
.data_in(VMR_L5D3_VMS_L5D3PHI2X1n6),
.enable(VMR_L5D3_VMS_L5D3PHI2X1n6_wr_en),
.number_out(VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1_number),
.read_add(VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1_read_add),
.data_out(VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X2;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2_read_add;
wire [13:0] VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2;
VMProjections  VMPROJ_L1L2_L5D3PHI2X2(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X2),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X2_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2_number),
.read_add(VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2),
.start(PR_L5D3_L1L2_start),
.done(VMPROJ_L1L2_L5D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI2X2n6;
wire VMR_L5D3_VMS_L5D3PHI2X2n6_wr_en;
wire [5:0] VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2_number;
wire [10:0] VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2_read_add;
wire [18:0] VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2;
VMStubs #("Match") VMS_L5D3PHI2X2n6(
.data_in(VMR_L5D3_VMS_L5D3PHI2X2n6),
.enable(VMR_L5D3_VMS_L5D3PHI2X2n6_wr_en),
.number_out(VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2_number),
.read_add(VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2_read_add),
.data_out(VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X1;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1_read_add;
wire [13:0] VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1;
VMProjections  VMPROJ_L1L2_L5D3PHI3X1(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X1),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X1_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1_number),
.read_add(VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1),
.start(PR_L5D3_L1L2_start),
.done(VMPROJ_L1L2_L5D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X1n6;
wire VMR_L5D3_VMS_L5D3PHI3X1n6_wr_en;
wire [5:0] VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1_number;
wire [10:0] VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1_read_add;
wire [18:0] VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1;
VMStubs #("Match") VMS_L5D3PHI3X1n6(
.data_in(VMR_L5D3_VMS_L5D3PHI3X1n6),
.enable(VMR_L5D3_VMS_L5D3PHI3X1n6_wr_en),
.number_out(VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1_number),
.read_add(VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1_read_add),
.data_out(VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X2;
wire PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2_number;
wire [8:0] VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2_read_add;
wire [13:0] VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2;
VMProjections  VMPROJ_L1L2_L5D3PHI3X2(
.data_in(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X2),
.enable(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X2_wr_en),
.number_out(VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2_number),
.read_add(VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2_read_add),
.data_out(VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2),
.start(PR_L5D3_L1L2_start),
.done(VMPROJ_L1L2_L5D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D3_VMS_L5D3PHI3X2n6;
wire VMR_L5D3_VMS_L5D3PHI3X2n6_wr_en;
wire [5:0] VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2_number;
wire [10:0] VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2_read_add;
wire [18:0] VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2;
VMStubs #("Match") VMS_L5D3PHI3X2n6(
.data_in(VMR_L5D3_VMS_L5D3PHI3X2n6),
.enable(VMR_L5D3_VMS_L5D3PHI3X2n6_wr_en),
.number_out(VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2_number),
.read_add(VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2_read_add),
.data_out(VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2),
.start(VMR_L5D3_start),
.done(VMS_L5D3PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X1;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1_read_add;
wire [13:0] VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1;
VMProjections  VMPROJ_L1L2_L5D4PHI1X1(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X1),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X1_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1_number),
.read_add(VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1),
.start(PR_L5D4_L1L2_start),
.done(VMPROJ_L1L2_L5D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X1n6;
wire VMR_L5D4_VMS_L5D4PHI1X1n6_wr_en;
wire [5:0] VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1_number;
wire [10:0] VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1_read_add;
wire [18:0] VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1;
VMStubs #("Match") VMS_L5D4PHI1X1n6(
.data_in(VMR_L5D4_VMS_L5D4PHI1X1n6),
.enable(VMR_L5D4_VMS_L5D4PHI1X1n6_wr_en),
.number_out(VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1_number),
.read_add(VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1_read_add),
.data_out(VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X2;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2_read_add;
wire [13:0] VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2;
VMProjections  VMPROJ_L1L2_L5D4PHI1X2(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X2),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X2_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2_number),
.read_add(VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2),
.start(PR_L5D4_L1L2_start),
.done(VMPROJ_L1L2_L5D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI1X2n4;
wire VMR_L5D4_VMS_L5D4PHI1X2n4_wr_en;
wire [5:0] VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2_number;
wire [10:0] VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2_read_add;
wire [18:0] VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2;
VMStubs #("Match") VMS_L5D4PHI1X2n4(
.data_in(VMR_L5D4_VMS_L5D4PHI1X2n4),
.enable(VMR_L5D4_VMS_L5D4PHI1X2n4_wr_en),
.number_out(VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2_number),
.read_add(VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2_read_add),
.data_out(VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X1;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1_read_add;
wire [13:0] VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1;
VMProjections  VMPROJ_L1L2_L5D4PHI2X1(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X1),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X1_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1_number),
.read_add(VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1),
.start(PR_L5D4_L1L2_start),
.done(VMPROJ_L1L2_L5D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X1n6;
wire VMR_L5D4_VMS_L5D4PHI2X1n6_wr_en;
wire [5:0] VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1_number;
wire [10:0] VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1_read_add;
wire [18:0] VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1;
VMStubs #("Match") VMS_L5D4PHI2X1n6(
.data_in(VMR_L5D4_VMS_L5D4PHI2X1n6),
.enable(VMR_L5D4_VMS_L5D4PHI2X1n6_wr_en),
.number_out(VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1_number),
.read_add(VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1_read_add),
.data_out(VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X2;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2_read_add;
wire [13:0] VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2;
VMProjections  VMPROJ_L1L2_L5D4PHI2X2(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X2),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X2_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2_number),
.read_add(VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2),
.start(PR_L5D4_L1L2_start),
.done(VMPROJ_L1L2_L5D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI2X2n4;
wire VMR_L5D4_VMS_L5D4PHI2X2n4_wr_en;
wire [5:0] VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2_number;
wire [10:0] VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2_read_add;
wire [18:0] VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2;
VMStubs #("Match") VMS_L5D4PHI2X2n4(
.data_in(VMR_L5D4_VMS_L5D4PHI2X2n4),
.enable(VMR_L5D4_VMS_L5D4PHI2X2n4_wr_en),
.number_out(VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2_number),
.read_add(VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2_read_add),
.data_out(VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X1;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1_read_add;
wire [13:0] VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1;
VMProjections  VMPROJ_L1L2_L5D4PHI3X1(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X1),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X1_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1_number),
.read_add(VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1),
.start(PR_L5D4_L1L2_start),
.done(VMPROJ_L1L2_L5D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X1n6;
wire VMR_L5D4_VMS_L5D4PHI3X1n6_wr_en;
wire [5:0] VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1_number;
wire [10:0] VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1_read_add;
wire [18:0] VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1;
VMStubs #("Match") VMS_L5D4PHI3X1n6(
.data_in(VMR_L5D4_VMS_L5D4PHI3X1n6),
.enable(VMR_L5D4_VMS_L5D4PHI3X1n6_wr_en),
.number_out(VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1_number),
.read_add(VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1_read_add),
.data_out(VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X2;
wire PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2_number;
wire [8:0] VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2_read_add;
wire [13:0] VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2;
VMProjections  VMPROJ_L1L2_L5D4PHI3X2(
.data_in(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X2),
.enable(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X2_wr_en),
.number_out(VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2_number),
.read_add(VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2_read_add),
.data_out(VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2),
.start(PR_L5D4_L1L2_start),
.done(VMPROJ_L1L2_L5D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L5D4_VMS_L5D4PHI3X2n4;
wire VMR_L5D4_VMS_L5D4PHI3X2n4_wr_en;
wire [5:0] VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2_number;
wire [10:0] VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2_read_add;
wire [18:0] VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2;
VMStubs #("Match") VMS_L5D4PHI3X2n4(
.data_in(VMR_L5D4_VMS_L5D4PHI3X2n4),
.enable(VMR_L5D4_VMS_L5D4PHI3X2n4_wr_en),
.number_out(VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2_number),
.read_add(VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2_read_add),
.data_out(VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2),
.start(VMR_L5D4_start),
.done(VMS_L5D4PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X1;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1_read_add;
wire [13:0] VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1;
VMProjections  VMPROJ_L1L2_L6D3PHI1X1(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X1),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X1_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1_number),
.read_add(VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1),
.start(PR_L6D3_L1L2_start),
.done(VMPROJ_L1L2_L6D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI1X1n3;
wire VMR_L6D3_VMS_L6D3PHI1X1n3_wr_en;
wire [5:0] VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1_number;
wire [10:0] VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1_read_add;
wire [18:0] VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1;
VMStubs #("Match") VMS_L6D3PHI1X1n3(
.data_in(VMR_L6D3_VMS_L6D3PHI1X1n3),
.enable(VMR_L6D3_VMS_L6D3PHI1X1n3_wr_en),
.number_out(VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1_number),
.read_add(VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1_read_add),
.data_out(VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X2;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2_read_add;
wire [13:0] VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2;
VMProjections  VMPROJ_L1L2_L6D3PHI1X2(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X2),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X2_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2_number),
.read_add(VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2),
.start(PR_L6D3_L1L2_start),
.done(VMPROJ_L1L2_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI1X2n4;
wire VMR_L6D3_VMS_L6D3PHI1X2n4_wr_en;
wire [5:0] VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2_number;
wire [10:0] VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2_read_add;
wire [18:0] VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2;
VMStubs #("Match") VMS_L6D3PHI1X2n4(
.data_in(VMR_L6D3_VMS_L6D3PHI1X2n4),
.enable(VMR_L6D3_VMS_L6D3PHI1X2n4_wr_en),
.number_out(VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2_number),
.read_add(VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2_read_add),
.data_out(VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X1;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1_read_add;
wire [13:0] VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1;
VMProjections  VMPROJ_L1L2_L6D3PHI2X1(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X1),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X1_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1_number),
.read_add(VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1),
.start(PR_L6D3_L1L2_start),
.done(VMPROJ_L1L2_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X1n4;
wire VMR_L6D3_VMS_L6D3PHI2X1n4_wr_en;
wire [5:0] VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1_number;
wire [10:0] VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1_read_add;
wire [18:0] VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1;
VMStubs #("Match") VMS_L6D3PHI2X1n4(
.data_in(VMR_L6D3_VMS_L6D3PHI2X1n4),
.enable(VMR_L6D3_VMS_L6D3PHI2X1n4_wr_en),
.number_out(VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1_number),
.read_add(VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1_read_add),
.data_out(VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X2;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2_read_add;
wire [13:0] VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2;
VMProjections  VMPROJ_L1L2_L6D3PHI2X2(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X2),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X2_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2_number),
.read_add(VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2),
.start(PR_L6D3_L1L2_start),
.done(VMPROJ_L1L2_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI2X2n6;
wire VMR_L6D3_VMS_L6D3PHI2X2n6_wr_en;
wire [5:0] VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2_number;
wire [10:0] VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2_read_add;
wire [18:0] VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2;
VMStubs #("Match") VMS_L6D3PHI2X2n6(
.data_in(VMR_L6D3_VMS_L6D3PHI2X2n6),
.enable(VMR_L6D3_VMS_L6D3PHI2X2n6_wr_en),
.number_out(VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2_number),
.read_add(VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2_read_add),
.data_out(VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X1;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1_read_add;
wire [13:0] VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1;
VMProjections  VMPROJ_L1L2_L6D3PHI3X1(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X1),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X1_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1_number),
.read_add(VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1),
.start(PR_L6D3_L1L2_start),
.done(VMPROJ_L1L2_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X1n4;
wire VMR_L6D3_VMS_L6D3PHI3X1n4_wr_en;
wire [5:0] VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1_number;
wire [10:0] VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1_read_add;
wire [18:0] VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1;
VMStubs #("Match") VMS_L6D3PHI3X1n4(
.data_in(VMR_L6D3_VMS_L6D3PHI3X1n4),
.enable(VMR_L6D3_VMS_L6D3PHI3X1n4_wr_en),
.number_out(VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1_number),
.read_add(VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1_read_add),
.data_out(VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X2;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2_read_add;
wire [13:0] VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2;
VMProjections  VMPROJ_L1L2_L6D3PHI3X2(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X2),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X2_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2_number),
.read_add(VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2),
.start(PR_L6D3_L1L2_start),
.done(VMPROJ_L1L2_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI3X2n6;
wire VMR_L6D3_VMS_L6D3PHI3X2n6_wr_en;
wire [5:0] VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2_number;
wire [10:0] VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2_read_add;
wire [18:0] VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2;
VMStubs #("Match") VMS_L6D3PHI3X2n6(
.data_in(VMR_L6D3_VMS_L6D3PHI3X2n6),
.enable(VMR_L6D3_VMS_L6D3PHI3X2n6_wr_en),
.number_out(VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2_number),
.read_add(VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2_read_add),
.data_out(VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X1;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1_read_add;
wire [13:0] VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1;
VMProjections  VMPROJ_L1L2_L6D3PHI4X1(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X1),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X1_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1_number),
.read_add(VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1),
.start(PR_L6D3_L1L2_start),
.done(VMPROJ_L1L2_L6D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI4X1n3;
wire VMR_L6D3_VMS_L6D3PHI4X1n3_wr_en;
wire [5:0] VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1_number;
wire [10:0] VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1_read_add;
wire [18:0] VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1;
VMStubs #("Match") VMS_L6D3PHI4X1n3(
.data_in(VMR_L6D3_VMS_L6D3PHI4X1n3),
.enable(VMR_L6D3_VMS_L6D3PHI4X1n3_wr_en),
.number_out(VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1_number),
.read_add(VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1_read_add),
.data_out(VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI4X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X2;
wire PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2_number;
wire [8:0] VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2_read_add;
wire [13:0] VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2;
VMProjections  VMPROJ_L1L2_L6D3PHI4X2(
.data_in(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X2),
.enable(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X2_wr_en),
.number_out(VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2_number),
.read_add(VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2_read_add),
.data_out(VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2),
.start(PR_L6D3_L1L2_start),
.done(VMPROJ_L1L2_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D3_VMS_L6D3PHI4X2n4;
wire VMR_L6D3_VMS_L6D3PHI4X2n4_wr_en;
wire [5:0] VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2_number;
wire [10:0] VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2_read_add;
wire [18:0] VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2;
VMStubs #("Match") VMS_L6D3PHI4X2n4(
.data_in(VMR_L6D3_VMS_L6D3PHI4X2n4),
.enable(VMR_L6D3_VMS_L6D3PHI4X2n4_wr_en),
.number_out(VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2_number),
.read_add(VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2_read_add),
.data_out(VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2),
.start(VMR_L6D3_start),
.done(VMS_L6D3PHI4X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X1;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1_read_add;
wire [13:0] VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1;
VMProjections  VMPROJ_L1L2_L6D4PHI1X1(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X1),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X1_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1_number),
.read_add(VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1),
.start(PR_L6D4_L1L2_start),
.done(VMPROJ_L1L2_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI1X1n4;
wire VMR_L6D4_VMS_L6D4PHI1X1n4_wr_en;
wire [5:0] VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1_number;
wire [10:0] VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1_read_add;
wire [18:0] VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1;
VMStubs #("Match") VMS_L6D4PHI1X1n4(
.data_in(VMR_L6D4_VMS_L6D4PHI1X1n4),
.enable(VMR_L6D4_VMS_L6D4PHI1X1n4_wr_en),
.number_out(VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1_number),
.read_add(VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1_read_add),
.data_out(VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X2;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2_read_add;
wire [13:0] VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2;
VMProjections  VMPROJ_L1L2_L6D4PHI1X2(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X2),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X2_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2_number),
.read_add(VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2),
.start(PR_L6D4_L1L2_start),
.done(VMPROJ_L1L2_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI1X2n4;
wire VMR_L6D4_VMS_L6D4PHI1X2n4_wr_en;
wire [5:0] VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2_number;
wire [10:0] VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2_read_add;
wire [18:0] VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2;
VMStubs #("Match") VMS_L6D4PHI1X2n4(
.data_in(VMR_L6D4_VMS_L6D4PHI1X2n4),
.enable(VMR_L6D4_VMS_L6D4PHI1X2n4_wr_en),
.number_out(VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2_number),
.read_add(VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2_read_add),
.data_out(VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X1;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1_read_add;
wire [13:0] VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1;
VMProjections  VMPROJ_L1L2_L6D4PHI2X1(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X1),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X1_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1_number),
.read_add(VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1),
.start(PR_L6D4_L1L2_start),
.done(VMPROJ_L1L2_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X1n6;
wire VMR_L6D4_VMS_L6D4PHI2X1n6_wr_en;
wire [5:0] VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1_number;
wire [10:0] VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1_read_add;
wire [18:0] VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1;
VMStubs #("Match") VMS_L6D4PHI2X1n6(
.data_in(VMR_L6D4_VMS_L6D4PHI2X1n6),
.enable(VMR_L6D4_VMS_L6D4PHI2X1n6_wr_en),
.number_out(VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1_number),
.read_add(VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1_read_add),
.data_out(VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X2;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2_read_add;
wire [13:0] VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2;
VMProjections  VMPROJ_L1L2_L6D4PHI2X2(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X2),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X2_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2_number),
.read_add(VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2),
.start(PR_L6D4_L1L2_start),
.done(VMPROJ_L1L2_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI2X2n6;
wire VMR_L6D4_VMS_L6D4PHI2X2n6_wr_en;
wire [5:0] VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2_number;
wire [10:0] VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2_read_add;
wire [18:0] VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2;
VMStubs #("Match") VMS_L6D4PHI2X2n6(
.data_in(VMR_L6D4_VMS_L6D4PHI2X2n6),
.enable(VMR_L6D4_VMS_L6D4PHI2X2n6_wr_en),
.number_out(VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2_number),
.read_add(VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2_read_add),
.data_out(VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X1;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1_read_add;
wire [13:0] VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1;
VMProjections  VMPROJ_L1L2_L6D4PHI3X1(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X1),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X1_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1_number),
.read_add(VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1),
.start(PR_L6D4_L1L2_start),
.done(VMPROJ_L1L2_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X1n6;
wire VMR_L6D4_VMS_L6D4PHI3X1n6_wr_en;
wire [5:0] VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1_number;
wire [10:0] VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1_read_add;
wire [18:0] VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1;
VMStubs #("Match") VMS_L6D4PHI3X1n6(
.data_in(VMR_L6D4_VMS_L6D4PHI3X1n6),
.enable(VMR_L6D4_VMS_L6D4PHI3X1n6_wr_en),
.number_out(VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1_number),
.read_add(VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1_read_add),
.data_out(VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X2;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2_read_add;
wire [13:0] VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2;
VMProjections  VMPROJ_L1L2_L6D4PHI3X2(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X2),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X2_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2_number),
.read_add(VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2),
.start(PR_L6D4_L1L2_start),
.done(VMPROJ_L1L2_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI3X2n6;
wire VMR_L6D4_VMS_L6D4PHI3X2n6_wr_en;
wire [5:0] VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2_number;
wire [10:0] VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2_read_add;
wire [18:0] VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2;
VMStubs #("Match") VMS_L6D4PHI3X2n6(
.data_in(VMR_L6D4_VMS_L6D4PHI3X2n6),
.enable(VMR_L6D4_VMS_L6D4PHI3X2n6_wr_en),
.number_out(VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2_number),
.read_add(VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2_read_add),
.data_out(VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X1;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X1_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1_read_add;
wire [13:0] VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1;
VMProjections  VMPROJ_L1L2_L6D4PHI4X1(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X1),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X1_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1_number),
.read_add(VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1),
.start(PR_L6D4_L1L2_start),
.done(VMPROJ_L1L2_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI4X1n4;
wire VMR_L6D4_VMS_L6D4PHI4X1n4_wr_en;
wire [5:0] VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1_number;
wire [10:0] VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1_read_add;
wire [18:0] VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1;
VMStubs #("Match") VMS_L6D4PHI4X1n4(
.data_in(VMR_L6D4_VMS_L6D4PHI4X1n4),
.enable(VMR_L6D4_VMS_L6D4PHI4X1n4_wr_en),
.number_out(VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1_number),
.read_add(VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1_read_add),
.data_out(VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI4X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X2;
wire PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X2_wr_en;
wire [5:0] VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2_number;
wire [8:0] VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2_read_add;
wire [13:0] VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2;
VMProjections  VMPROJ_L1L2_L6D4PHI4X2(
.data_in(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X2),
.enable(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X2_wr_en),
.number_out(VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2_number),
.read_add(VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2_read_add),
.data_out(VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2),
.start(PR_L6D4_L1L2_start),
.done(VMPROJ_L1L2_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L6D4_VMS_L6D4PHI4X2n4;
wire VMR_L6D4_VMS_L6D4PHI4X2n4_wr_en;
wire [5:0] VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2_number;
wire [10:0] VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2_read_add;
wire [18:0] VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2;
VMStubs #("Match") VMS_L6D4PHI4X2n4(
.data_in(VMR_L6D4_VMS_L6D4PHI4X2n4),
.enable(VMR_L6D4_VMS_L6D4PHI4X2n4_wr_en),
.number_out(VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2_number),
.read_add(VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2_read_add),
.data_out(VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2),
.start(VMR_L6D4_start),
.done(VMS_L6D4PHI4X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X1;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1_read_add;
wire [13:0] VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1;
VMProjections  VMPROJ_L5L6_L1D3PHI1X1(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X1),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X1_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1_number),
.read_add(VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1),
.start(PR_L1D3_L5L6_start),
.done(VMPROJ_L5L6_L1D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X1n8;
wire VMR_L1D3_VMS_L1D3PHI1X1n8_wr_en;
wire [5:0] VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1_number;
wire [10:0] VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1_read_add;
wire [18:0] VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1;
VMStubs #("Match") VMS_L1D3PHI1X1n8(
.data_in(VMR_L1D3_VMS_L1D3PHI1X1n8),
.enable(VMR_L1D3_VMS_L1D3PHI1X1n8_wr_en),
.number_out(VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1_number),
.read_add(VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1_read_add),
.data_out(VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X1n8_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X2;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2_read_add;
wire [13:0] VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2;
VMProjections  VMPROJ_L5L6_L1D3PHI1X2(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X2),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X2_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2_number),
.read_add(VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2),
.start(PR_L1D3_L5L6_start),
.done(VMPROJ_L5L6_L1D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI1X2n8;
wire VMR_L1D3_VMS_L1D3PHI1X2n8_wr_en;
wire [5:0] VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2_number;
wire [10:0] VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2_read_add;
wire [18:0] VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2;
VMStubs #("Match") VMS_L1D3PHI1X2n8(
.data_in(VMR_L1D3_VMS_L1D3PHI1X2n8),
.enable(VMR_L1D3_VMS_L1D3PHI1X2n8_wr_en),
.number_out(VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2_number),
.read_add(VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2_read_add),
.data_out(VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI1X2n8_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X1;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1_read_add;
wire [13:0] VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1;
VMProjections  VMPROJ_L5L6_L1D3PHI2X1(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X1),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X1_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1_number),
.read_add(VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1),
.start(PR_L1D3_L5L6_start),
.done(VMPROJ_L5L6_L1D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X1n8;
wire VMR_L1D3_VMS_L1D3PHI2X1n8_wr_en;
wire [5:0] VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1_number;
wire [10:0] VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1_read_add;
wire [18:0] VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1;
VMStubs #("Match") VMS_L1D3PHI2X1n8(
.data_in(VMR_L1D3_VMS_L1D3PHI2X1n8),
.enable(VMR_L1D3_VMS_L1D3PHI2X1n8_wr_en),
.number_out(VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1_number),
.read_add(VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1_read_add),
.data_out(VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X1n8_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X2;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2_read_add;
wire [13:0] VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2;
VMProjections  VMPROJ_L5L6_L1D3PHI2X2(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X2),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X2_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2_number),
.read_add(VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2),
.start(PR_L1D3_L5L6_start),
.done(VMPROJ_L5L6_L1D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI2X2n8;
wire VMR_L1D3_VMS_L1D3PHI2X2n8_wr_en;
wire [5:0] VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2_number;
wire [10:0] VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2_read_add;
wire [18:0] VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2;
VMStubs #("Match") VMS_L1D3PHI2X2n8(
.data_in(VMR_L1D3_VMS_L1D3PHI2X2n8),
.enable(VMR_L1D3_VMS_L1D3PHI2X2n8_wr_en),
.number_out(VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2_number),
.read_add(VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2_read_add),
.data_out(VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI2X2n8_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X1;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1_read_add;
wire [13:0] VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1;
VMProjections  VMPROJ_L5L6_L1D3PHI3X1(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X1),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X1_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1_number),
.read_add(VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1),
.start(PR_L1D3_L5L6_start),
.done(VMPROJ_L5L6_L1D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X1n8;
wire VMR_L1D3_VMS_L1D3PHI3X1n8_wr_en;
wire [5:0] VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1_number;
wire [10:0] VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1_read_add;
wire [18:0] VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1;
VMStubs #("Match") VMS_L1D3PHI3X1n8(
.data_in(VMR_L1D3_VMS_L1D3PHI3X1n8),
.enable(VMR_L1D3_VMS_L1D3PHI3X1n8_wr_en),
.number_out(VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1_number),
.read_add(VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1_read_add),
.data_out(VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X1n8_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X2;
wire PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2_number;
wire [8:0] VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2_read_add;
wire [13:0] VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2;
VMProjections  VMPROJ_L5L6_L1D3PHI3X2(
.data_in(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X2),
.enable(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X2_wr_en),
.number_out(VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2_number),
.read_add(VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2_read_add),
.data_out(VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2),
.start(PR_L1D3_L5L6_start),
.done(VMPROJ_L5L6_L1D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D3_VMS_L1D3PHI3X2n8;
wire VMR_L1D3_VMS_L1D3PHI3X2n8_wr_en;
wire [5:0] VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2_number;
wire [10:0] VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2_read_add;
wire [18:0] VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2;
VMStubs #("Match") VMS_L1D3PHI3X2n8(
.data_in(VMR_L1D3_VMS_L1D3PHI3X2n8),
.enable(VMR_L1D3_VMS_L1D3PHI3X2n8_wr_en),
.number_out(VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2_number),
.read_add(VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2_read_add),
.data_out(VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2),
.start(VMR_L1D3_start),
.done(VMS_L1D3PHI3X2n8_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X1;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1_read_add;
wire [13:0] VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1;
VMProjections  VMPROJ_L5L6_L1D4PHI1X1(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X1),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X1_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1_number),
.read_add(VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1),
.start(PR_L1D4_L5L6_start),
.done(VMPROJ_L5L6_L1D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI1X1n4;
wire VMR_L1D4_VMS_L1D4PHI1X1n4_wr_en;
wire [5:0] VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1_number;
wire [10:0] VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1_read_add;
wire [18:0] VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1;
VMStubs #("Match") VMS_L1D4PHI1X1n4(
.data_in(VMR_L1D4_VMS_L1D4PHI1X1n4),
.enable(VMR_L1D4_VMS_L1D4PHI1X1n4_wr_en),
.number_out(VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1_number),
.read_add(VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1_read_add),
.data_out(VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X2;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2_read_add;
wire [13:0] VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2;
VMProjections  VMPROJ_L5L6_L1D4PHI1X2(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X2),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X2_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2_number),
.read_add(VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2),
.start(PR_L1D4_L5L6_start),
.done(VMPROJ_L5L6_L1D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI1X2n2;
wire VMR_L1D4_VMS_L1D4PHI1X2n2_wr_en;
wire [5:0] VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2_number;
wire [10:0] VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2_read_add;
wire [18:0] VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2;
VMStubs #("Match") VMS_L1D4PHI1X2n2(
.data_in(VMR_L1D4_VMS_L1D4PHI1X2n2),
.enable(VMR_L1D4_VMS_L1D4PHI1X2n2_wr_en),
.number_out(VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2_number),
.read_add(VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2_read_add),
.data_out(VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI1X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X1;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1_read_add;
wire [13:0] VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1;
VMProjections  VMPROJ_L5L6_L1D4PHI2X1(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X1),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X1_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1_number),
.read_add(VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1),
.start(PR_L1D4_L5L6_start),
.done(VMPROJ_L5L6_L1D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI2X1n4;
wire VMR_L1D4_VMS_L1D4PHI2X1n4_wr_en;
wire [5:0] VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1_number;
wire [10:0] VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1_read_add;
wire [18:0] VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1;
VMStubs #("Match") VMS_L1D4PHI2X1n4(
.data_in(VMR_L1D4_VMS_L1D4PHI2X1n4),
.enable(VMR_L1D4_VMS_L1D4PHI2X1n4_wr_en),
.number_out(VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1_number),
.read_add(VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1_read_add),
.data_out(VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X2;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2_read_add;
wire [13:0] VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2;
VMProjections  VMPROJ_L5L6_L1D4PHI2X2(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X2),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X2_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2_number),
.read_add(VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2),
.start(PR_L1D4_L5L6_start),
.done(VMPROJ_L5L6_L1D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI2X2n2;
wire VMR_L1D4_VMS_L1D4PHI2X2n2_wr_en;
wire [5:0] VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2_number;
wire [10:0] VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2_read_add;
wire [18:0] VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2;
VMStubs #("Match") VMS_L1D4PHI2X2n2(
.data_in(VMR_L1D4_VMS_L1D4PHI2X2n2),
.enable(VMR_L1D4_VMS_L1D4PHI2X2n2_wr_en),
.number_out(VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2_number),
.read_add(VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2_read_add),
.data_out(VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI2X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X1;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1_read_add;
wire [13:0] VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1;
VMProjections  VMPROJ_L5L6_L1D4PHI3X1(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X1),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X1_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1_number),
.read_add(VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1),
.start(PR_L1D4_L5L6_start),
.done(VMPROJ_L5L6_L1D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI3X1n4;
wire VMR_L1D4_VMS_L1D4PHI3X1n4_wr_en;
wire [5:0] VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1_number;
wire [10:0] VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1_read_add;
wire [18:0] VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1;
VMStubs #("Match") VMS_L1D4PHI3X1n4(
.data_in(VMR_L1D4_VMS_L1D4PHI3X1n4),
.enable(VMR_L1D4_VMS_L1D4PHI3X1n4_wr_en),
.number_out(VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1_number),
.read_add(VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1_read_add),
.data_out(VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X2;
wire PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2_number;
wire [8:0] VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2_read_add;
wire [13:0] VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2;
VMProjections  VMPROJ_L5L6_L1D4PHI3X2(
.data_in(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X2),
.enable(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X2_wr_en),
.number_out(VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2_number),
.read_add(VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2_read_add),
.data_out(VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2),
.start(PR_L1D4_L5L6_start),
.done(VMPROJ_L5L6_L1D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L1D4_VMS_L1D4PHI3X2n2;
wire VMR_L1D4_VMS_L1D4PHI3X2n2_wr_en;
wire [5:0] VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2_number;
wire [10:0] VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2_read_add;
wire [18:0] VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2;
VMStubs #("Match") VMS_L1D4PHI3X2n2(
.data_in(VMR_L1D4_VMS_L1D4PHI3X2n2),
.enable(VMR_L1D4_VMS_L1D4PHI3X2n2_wr_en),
.number_out(VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2_number),
.read_add(VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2_read_add),
.data_out(VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2),
.start(VMR_L1D4_start),
.done(VMS_L1D4PHI3X2n2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X1;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1_read_add;
wire [13:0] VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1;
VMProjections  VMPROJ_L5L6_L2D3PHI1X1(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X1),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X1_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1_number),
.read_add(VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1),
.start(PR_L2D3_L5L6_start),
.done(VMPROJ_L5L6_L2D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI1X1n3;
wire VMR_L2D3_VMS_L2D3PHI1X1n3_wr_en;
wire [5:0] VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1_number;
wire [10:0] VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1_read_add;
wire [18:0] VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1;
VMStubs #("Match") VMS_L2D3PHI1X1n3(
.data_in(VMR_L2D3_VMS_L2D3PHI1X1n3),
.enable(VMR_L2D3_VMS_L2D3PHI1X1n3_wr_en),
.number_out(VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1_number),
.read_add(VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1_read_add),
.data_out(VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X2;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2_read_add;
wire [13:0] VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2;
VMProjections  VMPROJ_L5L6_L2D3PHI1X2(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X2),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X2_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2_number),
.read_add(VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2),
.start(PR_L2D3_L5L6_start),
.done(VMPROJ_L5L6_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI1X2n4;
wire VMR_L2D3_VMS_L2D3PHI1X2n4_wr_en;
wire [5:0] VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2_number;
wire [10:0] VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2_read_add;
wire [18:0] VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2;
VMStubs #("Match") VMS_L2D3PHI1X2n4(
.data_in(VMR_L2D3_VMS_L2D3PHI1X2n4),
.enable(VMR_L2D3_VMS_L2D3PHI1X2n4_wr_en),
.number_out(VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2_number),
.read_add(VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2_read_add),
.data_out(VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X1;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1_read_add;
wire [13:0] VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1;
VMProjections  VMPROJ_L5L6_L2D3PHI2X1(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X1),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X1_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1_number),
.read_add(VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1),
.start(PR_L2D3_L5L6_start),
.done(VMPROJ_L5L6_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X1n4;
wire VMR_L2D3_VMS_L2D3PHI2X1n4_wr_en;
wire [5:0] VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1_number;
wire [10:0] VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1_read_add;
wire [18:0] VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1;
VMStubs #("Match") VMS_L2D3PHI2X1n4(
.data_in(VMR_L2D3_VMS_L2D3PHI2X1n4),
.enable(VMR_L2D3_VMS_L2D3PHI2X1n4_wr_en),
.number_out(VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1_number),
.read_add(VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1_read_add),
.data_out(VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X2;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2_read_add;
wire [13:0] VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2;
VMProjections  VMPROJ_L5L6_L2D3PHI2X2(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X2),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X2_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2_number),
.read_add(VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2),
.start(PR_L2D3_L5L6_start),
.done(VMPROJ_L5L6_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI2X2n6;
wire VMR_L2D3_VMS_L2D3PHI2X2n6_wr_en;
wire [5:0] VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2_number;
wire [10:0] VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2_read_add;
wire [18:0] VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2;
VMStubs #("Match") VMS_L2D3PHI2X2n6(
.data_in(VMR_L2D3_VMS_L2D3PHI2X2n6),
.enable(VMR_L2D3_VMS_L2D3PHI2X2n6_wr_en),
.number_out(VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2_number),
.read_add(VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2_read_add),
.data_out(VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X1;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1_read_add;
wire [13:0] VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1;
VMProjections  VMPROJ_L5L6_L2D3PHI3X1(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X1),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X1_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1_number),
.read_add(VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1),
.start(PR_L2D3_L5L6_start),
.done(VMPROJ_L5L6_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X1n4;
wire VMR_L2D3_VMS_L2D3PHI3X1n4_wr_en;
wire [5:0] VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1_number;
wire [10:0] VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1_read_add;
wire [18:0] VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1;
VMStubs #("Match") VMS_L2D3PHI3X1n4(
.data_in(VMR_L2D3_VMS_L2D3PHI3X1n4),
.enable(VMR_L2D3_VMS_L2D3PHI3X1n4_wr_en),
.number_out(VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1_number),
.read_add(VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1_read_add),
.data_out(VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X2;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2_read_add;
wire [13:0] VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2;
VMProjections  VMPROJ_L5L6_L2D3PHI3X2(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X2),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X2_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2_number),
.read_add(VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2),
.start(PR_L2D3_L5L6_start),
.done(VMPROJ_L5L6_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI3X2n6;
wire VMR_L2D3_VMS_L2D3PHI3X2n6_wr_en;
wire [5:0] VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2_number;
wire [10:0] VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2_read_add;
wire [18:0] VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2;
VMStubs #("Match") VMS_L2D3PHI3X2n6(
.data_in(VMR_L2D3_VMS_L2D3PHI3X2n6),
.enable(VMR_L2D3_VMS_L2D3PHI3X2n6_wr_en),
.number_out(VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2_number),
.read_add(VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2_read_add),
.data_out(VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X1;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1_read_add;
wire [13:0] VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1;
VMProjections  VMPROJ_L5L6_L2D3PHI4X1(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X1),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X1_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1_number),
.read_add(VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1),
.start(PR_L2D3_L5L6_start),
.done(VMPROJ_L5L6_L2D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI4X1n3;
wire VMR_L2D3_VMS_L2D3PHI4X1n3_wr_en;
wire [5:0] VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1_number;
wire [10:0] VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1_read_add;
wire [18:0] VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1;
VMStubs #("Match") VMS_L2D3PHI4X1n3(
.data_in(VMR_L2D3_VMS_L2D3PHI4X1n3),
.enable(VMR_L2D3_VMS_L2D3PHI4X1n3_wr_en),
.number_out(VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1_number),
.read_add(VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1_read_add),
.data_out(VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI4X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X2;
wire PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2_number;
wire [8:0] VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2_read_add;
wire [13:0] VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2;
VMProjections  VMPROJ_L5L6_L2D3PHI4X2(
.data_in(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X2),
.enable(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X2_wr_en),
.number_out(VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2_number),
.read_add(VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2_read_add),
.data_out(VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2),
.start(PR_L2D3_L5L6_start),
.done(VMPROJ_L5L6_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D3_VMS_L2D3PHI4X2n4;
wire VMR_L2D3_VMS_L2D3PHI4X2n4_wr_en;
wire [5:0] VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2_number;
wire [10:0] VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2_read_add;
wire [18:0] VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2;
VMStubs #("Match") VMS_L2D3PHI4X2n4(
.data_in(VMR_L2D3_VMS_L2D3PHI4X2n4),
.enable(VMR_L2D3_VMS_L2D3PHI4X2n4_wr_en),
.number_out(VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2_number),
.read_add(VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2_read_add),
.data_out(VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2),
.start(VMR_L2D3_start),
.done(VMS_L2D3PHI4X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X1;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1_read_add;
wire [13:0] VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1;
VMProjections  VMPROJ_L5L6_L2D4PHI1X1(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X1),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X1_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1_number),
.read_add(VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1),
.start(PR_L2D4_L5L6_start),
.done(VMPROJ_L5L6_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI1X1n4;
wire VMR_L2D4_VMS_L2D4PHI1X1n4_wr_en;
wire [5:0] VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1_number;
wire [10:0] VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1_read_add;
wire [18:0] VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1;
VMStubs #("Match") VMS_L2D4PHI1X1n4(
.data_in(VMR_L2D4_VMS_L2D4PHI1X1n4),
.enable(VMR_L2D4_VMS_L2D4PHI1X1n4_wr_en),
.number_out(VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1_number),
.read_add(VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1_read_add),
.data_out(VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X2;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2_read_add;
wire [13:0] VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2;
VMProjections  VMPROJ_L5L6_L2D4PHI1X2(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X2),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X2_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2_number),
.read_add(VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2),
.start(PR_L2D4_L5L6_start),
.done(VMPROJ_L5L6_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI1X2n4;
wire VMR_L2D4_VMS_L2D4PHI1X2n4_wr_en;
wire [5:0] VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2_number;
wire [10:0] VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2_read_add;
wire [18:0] VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2;
VMStubs #("Match") VMS_L2D4PHI1X2n4(
.data_in(VMR_L2D4_VMS_L2D4PHI1X2n4),
.enable(VMR_L2D4_VMS_L2D4PHI1X2n4_wr_en),
.number_out(VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2_number),
.read_add(VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2_read_add),
.data_out(VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X1;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1_read_add;
wire [13:0] VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1;
VMProjections  VMPROJ_L5L6_L2D4PHI2X1(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X1),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X1_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1_number),
.read_add(VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1),
.start(PR_L2D4_L5L6_start),
.done(VMPROJ_L5L6_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X1n6;
wire VMR_L2D4_VMS_L2D4PHI2X1n6_wr_en;
wire [5:0] VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1_number;
wire [10:0] VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1_read_add;
wire [18:0] VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1;
VMStubs #("Match") VMS_L2D4PHI2X1n6(
.data_in(VMR_L2D4_VMS_L2D4PHI2X1n6),
.enable(VMR_L2D4_VMS_L2D4PHI2X1n6_wr_en),
.number_out(VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1_number),
.read_add(VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1_read_add),
.data_out(VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X2;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2_read_add;
wire [13:0] VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2;
VMProjections  VMPROJ_L5L6_L2D4PHI2X2(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X2),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X2_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2_number),
.read_add(VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2),
.start(PR_L2D4_L5L6_start),
.done(VMPROJ_L5L6_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI2X2n6;
wire VMR_L2D4_VMS_L2D4PHI2X2n6_wr_en;
wire [5:0] VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2_number;
wire [10:0] VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2_read_add;
wire [18:0] VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2;
VMStubs #("Match") VMS_L2D4PHI2X2n6(
.data_in(VMR_L2D4_VMS_L2D4PHI2X2n6),
.enable(VMR_L2D4_VMS_L2D4PHI2X2n6_wr_en),
.number_out(VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2_number),
.read_add(VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2_read_add),
.data_out(VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X1;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1_read_add;
wire [13:0] VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1;
VMProjections  VMPROJ_L5L6_L2D4PHI3X1(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X1),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X1_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1_number),
.read_add(VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1),
.start(PR_L2D4_L5L6_start),
.done(VMPROJ_L5L6_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X1n6;
wire VMR_L2D4_VMS_L2D4PHI3X1n6_wr_en;
wire [5:0] VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1_number;
wire [10:0] VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1_read_add;
wire [18:0] VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1;
VMStubs #("Match") VMS_L2D4PHI3X1n6(
.data_in(VMR_L2D4_VMS_L2D4PHI3X1n6),
.enable(VMR_L2D4_VMS_L2D4PHI3X1n6_wr_en),
.number_out(VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1_number),
.read_add(VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1_read_add),
.data_out(VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X2;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2_read_add;
wire [13:0] VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2;
VMProjections  VMPROJ_L5L6_L2D4PHI3X2(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X2),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X2_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2_number),
.read_add(VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2),
.start(PR_L2D4_L5L6_start),
.done(VMPROJ_L5L6_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI3X2n6;
wire VMR_L2D4_VMS_L2D4PHI3X2n6_wr_en;
wire [5:0] VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2_number;
wire [10:0] VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2_read_add;
wire [18:0] VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2;
VMStubs #("Match") VMS_L2D4PHI3X2n6(
.data_in(VMR_L2D4_VMS_L2D4PHI3X2n6),
.enable(VMR_L2D4_VMS_L2D4PHI3X2n6_wr_en),
.number_out(VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2_number),
.read_add(VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2_read_add),
.data_out(VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X1;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X1_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1_read_add;
wire [13:0] VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1;
VMProjections  VMPROJ_L5L6_L2D4PHI4X1(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X1),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X1_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1_number),
.read_add(VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1),
.start(PR_L2D4_L5L6_start),
.done(VMPROJ_L5L6_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI4X1n4;
wire VMR_L2D4_VMS_L2D4PHI4X1n4_wr_en;
wire [5:0] VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1_number;
wire [10:0] VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1_read_add;
wire [18:0] VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1;
VMStubs #("Match") VMS_L2D4PHI4X1n4(
.data_in(VMR_L2D4_VMS_L2D4PHI4X1n4),
.enable(VMR_L2D4_VMS_L2D4PHI4X1n4_wr_en),
.number_out(VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1_number),
.read_add(VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1_read_add),
.data_out(VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI4X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X2;
wire PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X2_wr_en;
wire [5:0] VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2_number;
wire [8:0] VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2_read_add;
wire [13:0] VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2;
VMProjections  VMPROJ_L5L6_L2D4PHI4X2(
.data_in(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X2),
.enable(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X2_wr_en),
.number_out(VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2_number),
.read_add(VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2_read_add),
.data_out(VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2),
.start(PR_L2D4_L5L6_start),
.done(VMPROJ_L5L6_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L2D4_VMS_L2D4PHI4X2n4;
wire VMR_L2D4_VMS_L2D4PHI4X2n4_wr_en;
wire [5:0] VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2_number;
wire [10:0] VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2_read_add;
wire [18:0] VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2;
VMStubs #("Match") VMS_L2D4PHI4X2n4(
.data_in(VMR_L2D4_VMS_L2D4PHI4X2n4),
.enable(VMR_L2D4_VMS_L2D4PHI4X2n4_wr_en),
.number_out(VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2_number),
.read_add(VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2_read_add),
.data_out(VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2),
.start(VMR_L2D4_start),
.done(VMS_L2D4PHI4X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X1;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1_read_add;
wire [13:0] VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1;
VMProjections  VMPROJ_L5L6_L3D3PHI1X1(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X1),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X1_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1_number),
.read_add(VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1),
.start(PR_L3D3_L5L6_start),
.done(VMPROJ_L5L6_L3D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X1n6;
wire VMR_L3D3_VMS_L3D3PHI1X1n6_wr_en;
wire [5:0] VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1_number;
wire [10:0] VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1_read_add;
wire [18:0] VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1;
VMStubs #("Match") VMS_L3D3PHI1X1n6(
.data_in(VMR_L3D3_VMS_L3D3PHI1X1n6),
.enable(VMR_L3D3_VMS_L3D3PHI1X1n6_wr_en),
.number_out(VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1_number),
.read_add(VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1_read_add),
.data_out(VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X2;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2_read_add;
wire [13:0] VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2;
VMProjections  VMPROJ_L5L6_L3D3PHI1X2(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X2),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X2_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2_number),
.read_add(VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2),
.start(PR_L3D3_L5L6_start),
.done(VMPROJ_L5L6_L3D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI1X2n6;
wire VMR_L3D3_VMS_L3D3PHI1X2n6_wr_en;
wire [5:0] VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2_number;
wire [10:0] VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2_read_add;
wire [18:0] VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2;
VMStubs #("Match") VMS_L3D3PHI1X2n6(
.data_in(VMR_L3D3_VMS_L3D3PHI1X2n6),
.enable(VMR_L3D3_VMS_L3D3PHI1X2n6_wr_en),
.number_out(VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2_number),
.read_add(VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2_read_add),
.data_out(VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI1X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X1;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1_read_add;
wire [13:0] VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1;
VMProjections  VMPROJ_L5L6_L3D3PHI2X1(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X1),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X1_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1_number),
.read_add(VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1),
.start(PR_L3D3_L5L6_start),
.done(VMPROJ_L5L6_L3D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X1n6;
wire VMR_L3D3_VMS_L3D3PHI2X1n6_wr_en;
wire [5:0] VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1_number;
wire [10:0] VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1_read_add;
wire [18:0] VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1;
VMStubs #("Match") VMS_L3D3PHI2X1n6(
.data_in(VMR_L3D3_VMS_L3D3PHI2X1n6),
.enable(VMR_L3D3_VMS_L3D3PHI2X1n6_wr_en),
.number_out(VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1_number),
.read_add(VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1_read_add),
.data_out(VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X2;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2_read_add;
wire [13:0] VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2;
VMProjections  VMPROJ_L5L6_L3D3PHI2X2(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X2),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X2_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2_number),
.read_add(VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2),
.start(PR_L3D3_L5L6_start),
.done(VMPROJ_L5L6_L3D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI2X2n6;
wire VMR_L3D3_VMS_L3D3PHI2X2n6_wr_en;
wire [5:0] VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2_number;
wire [10:0] VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2_read_add;
wire [18:0] VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2;
VMStubs #("Match") VMS_L3D3PHI2X2n6(
.data_in(VMR_L3D3_VMS_L3D3PHI2X2n6),
.enable(VMR_L3D3_VMS_L3D3PHI2X2n6_wr_en),
.number_out(VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2_number),
.read_add(VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2_read_add),
.data_out(VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X1;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1_read_add;
wire [13:0] VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1;
VMProjections  VMPROJ_L5L6_L3D3PHI3X1(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X1),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X1_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1_number),
.read_add(VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1),
.start(PR_L3D3_L5L6_start),
.done(VMPROJ_L5L6_L3D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X1n6;
wire VMR_L3D3_VMS_L3D3PHI3X1n6_wr_en;
wire [5:0] VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1_number;
wire [10:0] VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1_read_add;
wire [18:0] VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1;
VMStubs #("Match") VMS_L3D3PHI3X1n6(
.data_in(VMR_L3D3_VMS_L3D3PHI3X1n6),
.enable(VMR_L3D3_VMS_L3D3PHI3X1n6_wr_en),
.number_out(VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1_number),
.read_add(VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1_read_add),
.data_out(VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X2;
wire PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2_number;
wire [8:0] VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2_read_add;
wire [13:0] VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2;
VMProjections  VMPROJ_L5L6_L3D3PHI3X2(
.data_in(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X2),
.enable(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X2_wr_en),
.number_out(VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2_number),
.read_add(VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2_read_add),
.data_out(VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2),
.start(PR_L3D3_L5L6_start),
.done(VMPROJ_L5L6_L3D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D3_VMS_L3D3PHI3X2n6;
wire VMR_L3D3_VMS_L3D3PHI3X2n6_wr_en;
wire [5:0] VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2_number;
wire [10:0] VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2_read_add;
wire [18:0] VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2;
VMStubs #("Match") VMS_L3D3PHI3X2n6(
.data_in(VMR_L3D3_VMS_L3D3PHI3X2n6),
.enable(VMR_L3D3_VMS_L3D3PHI3X2n6_wr_en),
.number_out(VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2_number),
.read_add(VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2_read_add),
.data_out(VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2),
.start(VMR_L3D3_start),
.done(VMS_L3D3PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X1;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1_read_add;
wire [13:0] VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1;
VMProjections  VMPROJ_L5L6_L3D4PHI1X1(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X1),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X1_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1_number),
.read_add(VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1),
.start(PR_L3D4_L5L6_start),
.done(VMPROJ_L5L6_L3D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X1n6;
wire VMR_L3D4_VMS_L3D4PHI1X1n6_wr_en;
wire [5:0] VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1_number;
wire [10:0] VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1_read_add;
wire [18:0] VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1;
VMStubs #("Match") VMS_L3D4PHI1X1n6(
.data_in(VMR_L3D4_VMS_L3D4PHI1X1n6),
.enable(VMR_L3D4_VMS_L3D4PHI1X1n6_wr_en),
.number_out(VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1_number),
.read_add(VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1_read_add),
.data_out(VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X2;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2_read_add;
wire [13:0] VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2;
VMProjections  VMPROJ_L5L6_L3D4PHI1X2(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X2),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X2_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2_number),
.read_add(VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2),
.start(PR_L3D4_L5L6_start),
.done(VMPROJ_L5L6_L3D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI1X2n4;
wire VMR_L3D4_VMS_L3D4PHI1X2n4_wr_en;
wire [5:0] VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2_number;
wire [10:0] VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2_read_add;
wire [18:0] VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2;
VMStubs #("Match") VMS_L3D4PHI1X2n4(
.data_in(VMR_L3D4_VMS_L3D4PHI1X2n4),
.enable(VMR_L3D4_VMS_L3D4PHI1X2n4_wr_en),
.number_out(VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2_number),
.read_add(VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2_read_add),
.data_out(VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X1;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1_read_add;
wire [13:0] VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1;
VMProjections  VMPROJ_L5L6_L3D4PHI2X1(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X1),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X1_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1_number),
.read_add(VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1),
.start(PR_L3D4_L5L6_start),
.done(VMPROJ_L5L6_L3D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X1n6;
wire VMR_L3D4_VMS_L3D4PHI2X1n6_wr_en;
wire [5:0] VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1_number;
wire [10:0] VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1_read_add;
wire [18:0] VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1;
VMStubs #("Match") VMS_L3D4PHI2X1n6(
.data_in(VMR_L3D4_VMS_L3D4PHI2X1n6),
.enable(VMR_L3D4_VMS_L3D4PHI2X1n6_wr_en),
.number_out(VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1_number),
.read_add(VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1_read_add),
.data_out(VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X2;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2_read_add;
wire [13:0] VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2;
VMProjections  VMPROJ_L5L6_L3D4PHI2X2(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X2),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X2_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2_number),
.read_add(VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2),
.start(PR_L3D4_L5L6_start),
.done(VMPROJ_L5L6_L3D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI2X2n4;
wire VMR_L3D4_VMS_L3D4PHI2X2n4_wr_en;
wire [5:0] VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2_number;
wire [10:0] VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2_read_add;
wire [18:0] VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2;
VMStubs #("Match") VMS_L3D4PHI2X2n4(
.data_in(VMR_L3D4_VMS_L3D4PHI2X2n4),
.enable(VMR_L3D4_VMS_L3D4PHI2X2n4_wr_en),
.number_out(VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2_number),
.read_add(VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2_read_add),
.data_out(VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI2X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X1;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1_read_add;
wire [13:0] VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1;
VMProjections  VMPROJ_L5L6_L3D4PHI3X1(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X1),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X1_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1_number),
.read_add(VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1),
.start(PR_L3D4_L5L6_start),
.done(VMPROJ_L5L6_L3D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X1n6;
wire VMR_L3D4_VMS_L3D4PHI3X1n6_wr_en;
wire [5:0] VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1_number;
wire [10:0] VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1_read_add;
wire [18:0] VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1;
VMStubs #("Match") VMS_L3D4PHI3X1n6(
.data_in(VMR_L3D4_VMS_L3D4PHI3X1n6),
.enable(VMR_L3D4_VMS_L3D4PHI3X1n6_wr_en),
.number_out(VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1_number),
.read_add(VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1_read_add),
.data_out(VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X2;
wire PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2_number;
wire [8:0] VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2_read_add;
wire [13:0] VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2;
VMProjections  VMPROJ_L5L6_L3D4PHI3X2(
.data_in(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X2),
.enable(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X2_wr_en),
.number_out(VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2_number),
.read_add(VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2_read_add),
.data_out(VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2),
.start(PR_L3D4_L5L6_start),
.done(VMPROJ_L5L6_L3D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L3D4_VMS_L3D4PHI3X2n4;
wire VMR_L3D4_VMS_L3D4PHI3X2n4_wr_en;
wire [5:0] VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2_number;
wire [10:0] VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2_read_add;
wire [18:0] VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2;
VMStubs #("Match") VMS_L3D4PHI3X2n4(
.data_in(VMR_L3D4_VMS_L3D4PHI3X2n4),
.enable(VMR_L3D4_VMS_L3D4PHI3X2n4_wr_en),
.number_out(VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2_number),
.read_add(VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2_read_add),
.data_out(VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2),
.start(VMR_L3D4_start),
.done(VMS_L3D4PHI3X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X1;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1_read_add;
wire [13:0] VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1;
VMProjections  VMPROJ_L5L6_L4D3PHI1X1(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X1),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X1_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1_number),
.read_add(VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1),
.start(PR_L4D3_L5L6_start),
.done(VMPROJ_L5L6_L4D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI1X1n3;
wire VMR_L4D3_VMS_L4D3PHI1X1n3_wr_en;
wire [5:0] VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1_number;
wire [10:0] VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1_read_add;
wire [18:0] VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1;
VMStubs #("Match") VMS_L4D3PHI1X1n3(
.data_in(VMR_L4D3_VMS_L4D3PHI1X1n3),
.enable(VMR_L4D3_VMS_L4D3PHI1X1n3_wr_en),
.number_out(VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1_number),
.read_add(VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1_read_add),
.data_out(VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI1X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X2;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2_read_add;
wire [13:0] VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2;
VMProjections  VMPROJ_L5L6_L4D3PHI1X2(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X2),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X2_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2_number),
.read_add(VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2),
.start(PR_L4D3_L5L6_start),
.done(VMPROJ_L5L6_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI1X2n4;
wire VMR_L4D3_VMS_L4D3PHI1X2n4_wr_en;
wire [5:0] VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2_number;
wire [10:0] VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2_read_add;
wire [18:0] VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2;
VMStubs #("Match") VMS_L4D3PHI1X2n4(
.data_in(VMR_L4D3_VMS_L4D3PHI1X2n4),
.enable(VMR_L4D3_VMS_L4D3PHI1X2n4_wr_en),
.number_out(VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2_number),
.read_add(VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2_read_add),
.data_out(VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X1;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1_read_add;
wire [13:0] VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1;
VMProjections  VMPROJ_L5L6_L4D3PHI2X1(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X1),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X1_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1_number),
.read_add(VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1),
.start(PR_L4D3_L5L6_start),
.done(VMPROJ_L5L6_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X1n4;
wire VMR_L4D3_VMS_L4D3PHI2X1n4_wr_en;
wire [5:0] VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1_number;
wire [10:0] VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1_read_add;
wire [18:0] VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1;
VMStubs #("Match") VMS_L4D3PHI2X1n4(
.data_in(VMR_L4D3_VMS_L4D3PHI2X1n4),
.enable(VMR_L4D3_VMS_L4D3PHI2X1n4_wr_en),
.number_out(VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1_number),
.read_add(VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1_read_add),
.data_out(VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X2;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2_read_add;
wire [13:0] VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2;
VMProjections  VMPROJ_L5L6_L4D3PHI2X2(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X2),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X2_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2_number),
.read_add(VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2),
.start(PR_L4D3_L5L6_start),
.done(VMPROJ_L5L6_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI2X2n6;
wire VMR_L4D3_VMS_L4D3PHI2X2n6_wr_en;
wire [5:0] VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2_number;
wire [10:0] VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2_read_add;
wire [18:0] VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2;
VMStubs #("Match") VMS_L4D3PHI2X2n6(
.data_in(VMR_L4D3_VMS_L4D3PHI2X2n6),
.enable(VMR_L4D3_VMS_L4D3PHI2X2n6_wr_en),
.number_out(VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2_number),
.read_add(VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2_read_add),
.data_out(VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X1;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1_read_add;
wire [13:0] VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1;
VMProjections  VMPROJ_L5L6_L4D3PHI3X1(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X1),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X1_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1_number),
.read_add(VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1),
.start(PR_L4D3_L5L6_start),
.done(VMPROJ_L5L6_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X1n4;
wire VMR_L4D3_VMS_L4D3PHI3X1n4_wr_en;
wire [5:0] VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1_number;
wire [10:0] VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1_read_add;
wire [18:0] VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1;
VMStubs #("Match") VMS_L4D3PHI3X1n4(
.data_in(VMR_L4D3_VMS_L4D3PHI3X1n4),
.enable(VMR_L4D3_VMS_L4D3PHI3X1n4_wr_en),
.number_out(VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1_number),
.read_add(VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1_read_add),
.data_out(VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X2;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2_read_add;
wire [13:0] VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2;
VMProjections  VMPROJ_L5L6_L4D3PHI3X2(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X2),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X2_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2_number),
.read_add(VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2),
.start(PR_L4D3_L5L6_start),
.done(VMPROJ_L5L6_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI3X2n6;
wire VMR_L4D3_VMS_L4D3PHI3X2n6_wr_en;
wire [5:0] VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2_number;
wire [10:0] VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2_read_add;
wire [18:0] VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2;
VMStubs #("Match") VMS_L4D3PHI3X2n6(
.data_in(VMR_L4D3_VMS_L4D3PHI3X2n6),
.enable(VMR_L4D3_VMS_L4D3PHI3X2n6_wr_en),
.number_out(VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2_number),
.read_add(VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2_read_add),
.data_out(VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X1;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1_read_add;
wire [13:0] VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1;
VMProjections  VMPROJ_L5L6_L4D3PHI4X1(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X1),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X1_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1_number),
.read_add(VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1),
.start(PR_L4D3_L5L6_start),
.done(VMPROJ_L5L6_L4D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI4X1n3;
wire VMR_L4D3_VMS_L4D3PHI4X1n3_wr_en;
wire [5:0] VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1_number;
wire [10:0] VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1_read_add;
wire [18:0] VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1;
VMStubs #("Match") VMS_L4D3PHI4X1n3(
.data_in(VMR_L4D3_VMS_L4D3PHI4X1n3),
.enable(VMR_L4D3_VMS_L4D3PHI4X1n3_wr_en),
.number_out(VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1_number),
.read_add(VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1_read_add),
.data_out(VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI4X1n3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X2;
wire PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2_number;
wire [8:0] VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2_read_add;
wire [13:0] VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2;
VMProjections  VMPROJ_L5L6_L4D3PHI4X2(
.data_in(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X2),
.enable(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X2_wr_en),
.number_out(VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2_number),
.read_add(VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2_read_add),
.data_out(VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2),
.start(PR_L4D3_L5L6_start),
.done(VMPROJ_L5L6_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D3_VMS_L4D3PHI4X2n4;
wire VMR_L4D3_VMS_L4D3PHI4X2n4_wr_en;
wire [5:0] VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2_number;
wire [10:0] VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2_read_add;
wire [18:0] VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2;
VMStubs #("Match") VMS_L4D3PHI4X2n4(
.data_in(VMR_L4D3_VMS_L4D3PHI4X2n4),
.enable(VMR_L4D3_VMS_L4D3PHI4X2n4_wr_en),
.number_out(VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2_number),
.read_add(VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2_read_add),
.data_out(VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2),
.start(VMR_L4D3_start),
.done(VMS_L4D3PHI4X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X1;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1_read_add;
wire [13:0] VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1;
VMProjections  VMPROJ_L5L6_L4D4PHI1X1(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X1),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X1_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1_number),
.read_add(VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1),
.start(PR_L4D4_L5L6_start),
.done(VMPROJ_L5L6_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI1X1n4;
wire VMR_L4D4_VMS_L4D4PHI1X1n4_wr_en;
wire [5:0] VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1_number;
wire [10:0] VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1_read_add;
wire [18:0] VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1;
VMStubs #("Match") VMS_L4D4PHI1X1n4(
.data_in(VMR_L4D4_VMS_L4D4PHI1X1n4),
.enable(VMR_L4D4_VMS_L4D4PHI1X1n4_wr_en),
.number_out(VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1_number),
.read_add(VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1_read_add),
.data_out(VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI1X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X2;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2_read_add;
wire [13:0] VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2;
VMProjections  VMPROJ_L5L6_L4D4PHI1X2(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X2),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X2_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2_number),
.read_add(VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2),
.start(PR_L4D4_L5L6_start),
.done(VMPROJ_L5L6_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI1X2n4;
wire VMR_L4D4_VMS_L4D4PHI1X2n4_wr_en;
wire [5:0] VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2_number;
wire [10:0] VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2_read_add;
wire [18:0] VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2;
VMStubs #("Match") VMS_L4D4PHI1X2n4(
.data_in(VMR_L4D4_VMS_L4D4PHI1X2n4),
.enable(VMR_L4D4_VMS_L4D4PHI1X2n4_wr_en),
.number_out(VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2_number),
.read_add(VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2_read_add),
.data_out(VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI1X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X1;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1_read_add;
wire [13:0] VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1;
VMProjections  VMPROJ_L5L6_L4D4PHI2X1(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X1),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X1_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1_number),
.read_add(VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1),
.start(PR_L4D4_L5L6_start),
.done(VMPROJ_L5L6_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X1n6;
wire VMR_L4D4_VMS_L4D4PHI2X1n6_wr_en;
wire [5:0] VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1_number;
wire [10:0] VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1_read_add;
wire [18:0] VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1;
VMStubs #("Match") VMS_L4D4PHI2X1n6(
.data_in(VMR_L4D4_VMS_L4D4PHI2X1n6),
.enable(VMR_L4D4_VMS_L4D4PHI2X1n6_wr_en),
.number_out(VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1_number),
.read_add(VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1_read_add),
.data_out(VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X2;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2_read_add;
wire [13:0] VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2;
VMProjections  VMPROJ_L5L6_L4D4PHI2X2(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X2),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X2_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2_number),
.read_add(VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2),
.start(PR_L4D4_L5L6_start),
.done(VMPROJ_L5L6_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI2X2n6;
wire VMR_L4D4_VMS_L4D4PHI2X2n6_wr_en;
wire [5:0] VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2_number;
wire [10:0] VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2_read_add;
wire [18:0] VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2;
VMStubs #("Match") VMS_L4D4PHI2X2n6(
.data_in(VMR_L4D4_VMS_L4D4PHI2X2n6),
.enable(VMR_L4D4_VMS_L4D4PHI2X2n6_wr_en),
.number_out(VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2_number),
.read_add(VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2_read_add),
.data_out(VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI2X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X1;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1_read_add;
wire [13:0] VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1;
VMProjections  VMPROJ_L5L6_L4D4PHI3X1(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X1),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X1_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1_number),
.read_add(VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1),
.start(PR_L4D4_L5L6_start),
.done(VMPROJ_L5L6_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X1n6;
wire VMR_L4D4_VMS_L4D4PHI3X1n6_wr_en;
wire [5:0] VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1_number;
wire [10:0] VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1_read_add;
wire [18:0] VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1;
VMStubs #("Match") VMS_L4D4PHI3X1n6(
.data_in(VMR_L4D4_VMS_L4D4PHI3X1n6),
.enable(VMR_L4D4_VMS_L4D4PHI3X1n6_wr_en),
.number_out(VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1_number),
.read_add(VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1_read_add),
.data_out(VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X1n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X2;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2_read_add;
wire [13:0] VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2;
VMProjections  VMPROJ_L5L6_L4D4PHI3X2(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X2),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X2_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2_number),
.read_add(VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2),
.start(PR_L4D4_L5L6_start),
.done(VMPROJ_L5L6_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI3X2n6;
wire VMR_L4D4_VMS_L4D4PHI3X2n6_wr_en;
wire [5:0] VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2_number;
wire [10:0] VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2_read_add;
wire [18:0] VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2;
VMStubs #("Match") VMS_L4D4PHI3X2n6(
.data_in(VMR_L4D4_VMS_L4D4PHI3X2n6),
.enable(VMR_L4D4_VMS_L4D4PHI3X2n6_wr_en),
.number_out(VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2_number),
.read_add(VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2_read_add),
.data_out(VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI3X2n6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X1;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X1_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1_read_add;
wire [13:0] VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1;
VMProjections  VMPROJ_L5L6_L4D4PHI4X1(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X1),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X1_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1_number),
.read_add(VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1),
.start(PR_L4D4_L5L6_start),
.done(VMPROJ_L5L6_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI4X1n4;
wire VMR_L4D4_VMS_L4D4PHI4X1n4_wr_en;
wire [5:0] VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1_number;
wire [10:0] VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1_read_add;
wire [18:0] VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1;
VMStubs #("Match") VMS_L4D4PHI4X1n4(
.data_in(VMR_L4D4_VMS_L4D4PHI4X1n4),
.enable(VMR_L4D4_VMS_L4D4PHI4X1n4_wr_en),
.number_out(VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1_number),
.read_add(VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1_read_add),
.data_out(VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI4X1n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [13:0] PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X2;
wire PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X2_wr_en;
wire [5:0] VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2_number;
wire [8:0] VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2_read_add;
wire [13:0] VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2;
VMProjections  VMPROJ_L5L6_L4D4PHI4X2(
.data_in(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X2),
.enable(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X2_wr_en),
.number_out(VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2_number),
.read_add(VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2_read_add),
.data_out(VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2),
.start(PR_L4D4_L5L6_start),
.done(VMPROJ_L5L6_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [18:0] VMR_L4D4_VMS_L4D4PHI4X2n4;
wire VMR_L4D4_VMS_L4D4PHI4X2n4_wr_en;
wire [5:0] VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2_number;
wire [10:0] VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2_read_add;
wire [18:0] VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2;
VMStubs #("Match") VMS_L4D4PHI4X2n4(
.data_in(VMR_L4D4_VMS_L4D4PHI4X2n4),
.enable(VMR_L4D4_VMS_L4D4PHI4X2n4_wr_en),
.number_out(VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2_number),
.read_add(VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2_read_add),
.data_out(VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2),
.start(VMR_L4D4_start),
.done(VMS_L4D4PHI4X2n4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D3PHI1X1_CM_L3L4_L1D3PHI1X1;
wire ME_L3L4_L1D3PHI1X1_CM_L3L4_L1D3PHI1X1_wr_en;
wire [5:0] CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI1X1(
.data_in(ME_L3L4_L1D3PHI1X1_CM_L3L4_L1D3PHI1X1),
.enable(ME_L3L4_L1D3PHI1X1_CM_L3L4_L1D3PHI1X1_wr_en),
.number_out(CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3),
.start(ME_L3L4_L1D3PHI1X1_start),
.done(CM_L3L4_L1D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D3PHI1X2_CM_L3L4_L1D3PHI1X2;
wire ME_L3L4_L1D3PHI1X2_CM_L3L4_L1D3PHI1X2_wr_en;
wire [5:0] CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI1X2(
.data_in(ME_L3L4_L1D3PHI1X2_CM_L3L4_L1D3PHI1X2),
.enable(ME_L3L4_L1D3PHI1X2_CM_L3L4_L1D3PHI1X2_wr_en),
.number_out(CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3),
.start(ME_L3L4_L1D3PHI1X2_start),
.done(CM_L3L4_L1D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D3PHI2X1_CM_L3L4_L1D3PHI2X1;
wire ME_L3L4_L1D3PHI2X1_CM_L3L4_L1D3PHI2X1_wr_en;
wire [5:0] CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI2X1(
.data_in(ME_L3L4_L1D3PHI2X1_CM_L3L4_L1D3PHI2X1),
.enable(ME_L3L4_L1D3PHI2X1_CM_L3L4_L1D3PHI2X1_wr_en),
.number_out(CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3),
.start(ME_L3L4_L1D3PHI2X1_start),
.done(CM_L3L4_L1D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D3PHI2X2_CM_L3L4_L1D3PHI2X2;
wire ME_L3L4_L1D3PHI2X2_CM_L3L4_L1D3PHI2X2_wr_en;
wire [5:0] CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI2X2(
.data_in(ME_L3L4_L1D3PHI2X2_CM_L3L4_L1D3PHI2X2),
.enable(ME_L3L4_L1D3PHI2X2_CM_L3L4_L1D3PHI2X2_wr_en),
.number_out(CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3),
.start(ME_L3L4_L1D3PHI2X2_start),
.done(CM_L3L4_L1D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D3PHI3X1_CM_L3L4_L1D3PHI3X1;
wire ME_L3L4_L1D3PHI3X1_CM_L3L4_L1D3PHI3X1_wr_en;
wire [5:0] CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI3X1(
.data_in(ME_L3L4_L1D3PHI3X1_CM_L3L4_L1D3PHI3X1),
.enable(ME_L3L4_L1D3PHI3X1_CM_L3L4_L1D3PHI3X1_wr_en),
.number_out(CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3),
.start(ME_L3L4_L1D3PHI3X1_start),
.done(CM_L3L4_L1D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D3PHI3X2_CM_L3L4_L1D3PHI3X2;
wire ME_L3L4_L1D3PHI3X2_CM_L3L4_L1D3PHI3X2_wr_en;
wire [5:0] CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3_number;
wire [8:0] CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3_read_add;
wire [11:0] CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3;
CandidateMatch  CM_L3L4_L1D3PHI3X2(
.data_in(ME_L3L4_L1D3PHI3X2_CM_L3L4_L1D3PHI3X2),
.enable(ME_L3L4_L1D3PHI3X2_CM_L3L4_L1D3PHI3X2_wr_en),
.number_out(CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3_number),
.read_add(CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3_read_add),
.data_out(CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3),
.start(ME_L3L4_L1D3PHI3X2_start),
.done(CM_L3L4_L1D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L1D3_L3L4_AP_L3L4_L1D3;
wire PR_L1D3_L3L4_AP_L3L4_L1D3_wr_en;
wire [8:0] AP_L3L4_L1D3_MC_L3L4_L1D3_read_add;
wire [55:0] AP_L3L4_L1D3_MC_L3L4_L1D3;
AllProj  AP_L3L4_L1D3(
.data_in(PR_L1D3_L3L4_AP_L3L4_L1D3),
.enable(PR_L1D3_L3L4_AP_L3L4_L1D3_wr_en),
.read_add(AP_L3L4_L1D3_MC_L3L4_L1D3_read_add),
.data_out(AP_L3L4_L1D3_MC_L3L4_L1D3),
.start(PR_L1D3_L3L4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L1D3_AS_L1D3n3;
wire VMR_L1D3_AS_L1D3n3_wr_en;
wire [10:0] AS_L1D3n3_MC_L3L4_L1D3_read_add;
wire [35:0] AS_L1D3n3_MC_L3L4_L1D3;
AllStubs  AS_L1D3n3(
.data_in(VMR_L1D3_AS_L1D3n3),
.enable(VMR_L1D3_AS_L1D3n3_wr_en),
.read_add_MC(AS_L1D3n3_MC_L3L4_L1D3_read_add),
.data_out_MC(AS_L1D3n3_MC_L3L4_L1D3),
.start(VMR_L1D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D4PHI1X1_CM_L3L4_L1D4PHI1X1;
wire ME_L3L4_L1D4PHI1X1_CM_L3L4_L1D4PHI1X1_wr_en;
wire [5:0] CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI1X1(
.data_in(ME_L3L4_L1D4PHI1X1_CM_L3L4_L1D4PHI1X1),
.enable(ME_L3L4_L1D4PHI1X1_CM_L3L4_L1D4PHI1X1_wr_en),
.number_out(CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4),
.start(ME_L3L4_L1D4PHI1X1_start),
.done(CM_L3L4_L1D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D4PHI1X2_CM_L3L4_L1D4PHI1X2;
wire ME_L3L4_L1D4PHI1X2_CM_L3L4_L1D4PHI1X2_wr_en;
wire [5:0] CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI1X2(
.data_in(ME_L3L4_L1D4PHI1X2_CM_L3L4_L1D4PHI1X2),
.enable(ME_L3L4_L1D4PHI1X2_CM_L3L4_L1D4PHI1X2_wr_en),
.number_out(CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4),
.start(ME_L3L4_L1D4PHI1X2_start),
.done(CM_L3L4_L1D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D4PHI2X1_CM_L3L4_L1D4PHI2X1;
wire ME_L3L4_L1D4PHI2X1_CM_L3L4_L1D4PHI2X1_wr_en;
wire [5:0] CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI2X1(
.data_in(ME_L3L4_L1D4PHI2X1_CM_L3L4_L1D4PHI2X1),
.enable(ME_L3L4_L1D4PHI2X1_CM_L3L4_L1D4PHI2X1_wr_en),
.number_out(CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4),
.start(ME_L3L4_L1D4PHI2X1_start),
.done(CM_L3L4_L1D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D4PHI2X2_CM_L3L4_L1D4PHI2X2;
wire ME_L3L4_L1D4PHI2X2_CM_L3L4_L1D4PHI2X2_wr_en;
wire [5:0] CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI2X2(
.data_in(ME_L3L4_L1D4PHI2X2_CM_L3L4_L1D4PHI2X2),
.enable(ME_L3L4_L1D4PHI2X2_CM_L3L4_L1D4PHI2X2_wr_en),
.number_out(CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4),
.start(ME_L3L4_L1D4PHI2X2_start),
.done(CM_L3L4_L1D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D4PHI3X1_CM_L3L4_L1D4PHI3X1;
wire ME_L3L4_L1D4PHI3X1_CM_L3L4_L1D4PHI3X1_wr_en;
wire [5:0] CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI3X1(
.data_in(ME_L3L4_L1D4PHI3X1_CM_L3L4_L1D4PHI3X1),
.enable(ME_L3L4_L1D4PHI3X1_CM_L3L4_L1D4PHI3X1_wr_en),
.number_out(CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4),
.start(ME_L3L4_L1D4PHI3X1_start),
.done(CM_L3L4_L1D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L1D4PHI3X2_CM_L3L4_L1D4PHI3X2;
wire ME_L3L4_L1D4PHI3X2_CM_L3L4_L1D4PHI3X2_wr_en;
wire [5:0] CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4_number;
wire [8:0] CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4_read_add;
wire [11:0] CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4;
CandidateMatch  CM_L3L4_L1D4PHI3X2(
.data_in(ME_L3L4_L1D4PHI3X2_CM_L3L4_L1D4PHI3X2),
.enable(ME_L3L4_L1D4PHI3X2_CM_L3L4_L1D4PHI3X2_wr_en),
.number_out(CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4_number),
.read_add(CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4_read_add),
.data_out(CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4),
.start(ME_L3L4_L1D4PHI3X2_start),
.done(CM_L3L4_L1D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L1D4_L3L4_AP_L3L4_L1D4;
wire PR_L1D4_L3L4_AP_L3L4_L1D4_wr_en;
wire [8:0] AP_L3L4_L1D4_MC_L3L4_L1D4_read_add;
wire [55:0] AP_L3L4_L1D4_MC_L3L4_L1D4;
AllProj  AP_L3L4_L1D4(
.data_in(PR_L1D4_L3L4_AP_L3L4_L1D4),
.enable(PR_L1D4_L3L4_AP_L3L4_L1D4_wr_en),
.read_add(AP_L3L4_L1D4_MC_L3L4_L1D4_read_add),
.data_out(AP_L3L4_L1D4_MC_L3L4_L1D4),
.start(PR_L1D4_L3L4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L1D4_AS_L1D4n2;
wire VMR_L1D4_AS_L1D4n2_wr_en;
wire [10:0] AS_L1D4n2_MC_L3L4_L1D4_read_add;
wire [35:0] AS_L1D4n2_MC_L3L4_L1D4;
AllStubs  AS_L1D4n2(
.data_in(VMR_L1D4_AS_L1D4n2),
.enable(VMR_L1D4_AS_L1D4n2_wr_en),
.read_add_MC(AS_L1D4n2_MC_L3L4_L1D4_read_add),
.data_out_MC(AS_L1D4n2_MC_L3L4_L1D4),
.start(VMR_L1D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D3PHI1X1_CM_L3L4_L2D3PHI1X1;
wire ME_L3L4_L2D3PHI1X1_CM_L3L4_L2D3PHI1X1_wr_en;
wire [5:0] CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI1X1(
.data_in(ME_L3L4_L2D3PHI1X1_CM_L3L4_L2D3PHI1X1),
.enable(ME_L3L4_L2D3PHI1X1_CM_L3L4_L2D3PHI1X1_wr_en),
.number_out(CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3),
.start(ME_L3L4_L2D3PHI1X1_start),
.done(CM_L3L4_L2D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D3PHI1X2_CM_L3L4_L2D3PHI1X2;
wire ME_L3L4_L2D3PHI1X2_CM_L3L4_L2D3PHI1X2_wr_en;
wire [5:0] CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI1X2(
.data_in(ME_L3L4_L2D3PHI1X2_CM_L3L4_L2D3PHI1X2),
.enable(ME_L3L4_L2D3PHI1X2_CM_L3L4_L2D3PHI1X2_wr_en),
.number_out(CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3),
.start(ME_L3L4_L2D3PHI1X2_start),
.done(CM_L3L4_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D3PHI2X1_CM_L3L4_L2D3PHI2X1;
wire ME_L3L4_L2D3PHI2X1_CM_L3L4_L2D3PHI2X1_wr_en;
wire [5:0] CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI2X1(
.data_in(ME_L3L4_L2D3PHI2X1_CM_L3L4_L2D3PHI2X1),
.enable(ME_L3L4_L2D3PHI2X1_CM_L3L4_L2D3PHI2X1_wr_en),
.number_out(CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3),
.start(ME_L3L4_L2D3PHI2X1_start),
.done(CM_L3L4_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D3PHI2X2_CM_L3L4_L2D3PHI2X2;
wire ME_L3L4_L2D3PHI2X2_CM_L3L4_L2D3PHI2X2_wr_en;
wire [5:0] CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI2X2(
.data_in(ME_L3L4_L2D3PHI2X2_CM_L3L4_L2D3PHI2X2),
.enable(ME_L3L4_L2D3PHI2X2_CM_L3L4_L2D3PHI2X2_wr_en),
.number_out(CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3),
.start(ME_L3L4_L2D3PHI2X2_start),
.done(CM_L3L4_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D3PHI3X1_CM_L3L4_L2D3PHI3X1;
wire ME_L3L4_L2D3PHI3X1_CM_L3L4_L2D3PHI3X1_wr_en;
wire [5:0] CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI3X1(
.data_in(ME_L3L4_L2D3PHI3X1_CM_L3L4_L2D3PHI3X1),
.enable(ME_L3L4_L2D3PHI3X1_CM_L3L4_L2D3PHI3X1_wr_en),
.number_out(CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3),
.start(ME_L3L4_L2D3PHI3X1_start),
.done(CM_L3L4_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D3PHI3X2_CM_L3L4_L2D3PHI3X2;
wire ME_L3L4_L2D3PHI3X2_CM_L3L4_L2D3PHI3X2_wr_en;
wire [5:0] CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI3X2(
.data_in(ME_L3L4_L2D3PHI3X2_CM_L3L4_L2D3PHI3X2),
.enable(ME_L3L4_L2D3PHI3X2_CM_L3L4_L2D3PHI3X2_wr_en),
.number_out(CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3),
.start(ME_L3L4_L2D3PHI3X2_start),
.done(CM_L3L4_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D3PHI4X1_CM_L3L4_L2D3PHI4X1;
wire ME_L3L4_L2D3PHI4X1_CM_L3L4_L2D3PHI4X1_wr_en;
wire [5:0] CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI4X1(
.data_in(ME_L3L4_L2D3PHI4X1_CM_L3L4_L2D3PHI4X1),
.enable(ME_L3L4_L2D3PHI4X1_CM_L3L4_L2D3PHI4X1_wr_en),
.number_out(CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3),
.start(ME_L3L4_L2D3PHI4X1_start),
.done(CM_L3L4_L2D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D3PHI4X2_CM_L3L4_L2D3PHI4X2;
wire ME_L3L4_L2D3PHI4X2_CM_L3L4_L2D3PHI4X2_wr_en;
wire [5:0] CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3_number;
wire [8:0] CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3_read_add;
wire [11:0] CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3;
CandidateMatch  CM_L3L4_L2D3PHI4X2(
.data_in(ME_L3L4_L2D3PHI4X2_CM_L3L4_L2D3PHI4X2),
.enable(ME_L3L4_L2D3PHI4X2_CM_L3L4_L2D3PHI4X2_wr_en),
.number_out(CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3_number),
.read_add(CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3_read_add),
.data_out(CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3),
.start(ME_L3L4_L2D3PHI4X2_start),
.done(CM_L3L4_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L2D3_L3L4_AP_L3L4_L2D3;
wire PR_L2D3_L3L4_AP_L3L4_L2D3_wr_en;
wire [8:0] AP_L3L4_L2D3_MC_L3L4_L2D3_read_add;
wire [55:0] AP_L3L4_L2D3_MC_L3L4_L2D3;
AllProj  AP_L3L4_L2D3(
.data_in(PR_L2D3_L3L4_AP_L3L4_L2D3),
.enable(PR_L2D3_L3L4_AP_L3L4_L2D3_wr_en),
.read_add(AP_L3L4_L2D3_MC_L3L4_L2D3_read_add),
.data_out(AP_L3L4_L2D3_MC_L3L4_L2D3),
.start(PR_L2D3_L3L4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L2D3_AS_L2D3n2;
wire VMR_L2D3_AS_L2D3n2_wr_en;
wire [10:0] AS_L2D3n2_MC_L3L4_L2D3_read_add;
wire [35:0] AS_L2D3n2_MC_L3L4_L2D3;
AllStubs  AS_L2D3n2(
.data_in(VMR_L2D3_AS_L2D3n2),
.enable(VMR_L2D3_AS_L2D3n2_wr_en),
.read_add_MC(AS_L2D3n2_MC_L3L4_L2D3_read_add),
.data_out_MC(AS_L2D3n2_MC_L3L4_L2D3),
.start(VMR_L2D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D4PHI1X1_CM_L3L4_L2D4PHI1X1;
wire ME_L3L4_L2D4PHI1X1_CM_L3L4_L2D4PHI1X1_wr_en;
wire [5:0] CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI1X1(
.data_in(ME_L3L4_L2D4PHI1X1_CM_L3L4_L2D4PHI1X1),
.enable(ME_L3L4_L2D4PHI1X1_CM_L3L4_L2D4PHI1X1_wr_en),
.number_out(CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4),
.start(ME_L3L4_L2D4PHI1X1_start),
.done(CM_L3L4_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D4PHI1X2_CM_L3L4_L2D4PHI1X2;
wire ME_L3L4_L2D4PHI1X2_CM_L3L4_L2D4PHI1X2_wr_en;
wire [5:0] CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI1X2(
.data_in(ME_L3L4_L2D4PHI1X2_CM_L3L4_L2D4PHI1X2),
.enable(ME_L3L4_L2D4PHI1X2_CM_L3L4_L2D4PHI1X2_wr_en),
.number_out(CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4),
.start(ME_L3L4_L2D4PHI1X2_start),
.done(CM_L3L4_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D4PHI2X1_CM_L3L4_L2D4PHI2X1;
wire ME_L3L4_L2D4PHI2X1_CM_L3L4_L2D4PHI2X1_wr_en;
wire [5:0] CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI2X1(
.data_in(ME_L3L4_L2D4PHI2X1_CM_L3L4_L2D4PHI2X1),
.enable(ME_L3L4_L2D4PHI2X1_CM_L3L4_L2D4PHI2X1_wr_en),
.number_out(CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4),
.start(ME_L3L4_L2D4PHI2X1_start),
.done(CM_L3L4_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D4PHI2X2_CM_L3L4_L2D4PHI2X2;
wire ME_L3L4_L2D4PHI2X2_CM_L3L4_L2D4PHI2X2_wr_en;
wire [5:0] CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI2X2(
.data_in(ME_L3L4_L2D4PHI2X2_CM_L3L4_L2D4PHI2X2),
.enable(ME_L3L4_L2D4PHI2X2_CM_L3L4_L2D4PHI2X2_wr_en),
.number_out(CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4),
.start(ME_L3L4_L2D4PHI2X2_start),
.done(CM_L3L4_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D4PHI3X1_CM_L3L4_L2D4PHI3X1;
wire ME_L3L4_L2D4PHI3X1_CM_L3L4_L2D4PHI3X1_wr_en;
wire [5:0] CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI3X1(
.data_in(ME_L3L4_L2D4PHI3X1_CM_L3L4_L2D4PHI3X1),
.enable(ME_L3L4_L2D4PHI3X1_CM_L3L4_L2D4PHI3X1_wr_en),
.number_out(CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4),
.start(ME_L3L4_L2D4PHI3X1_start),
.done(CM_L3L4_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D4PHI3X2_CM_L3L4_L2D4PHI3X2;
wire ME_L3L4_L2D4PHI3X2_CM_L3L4_L2D4PHI3X2_wr_en;
wire [5:0] CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI3X2(
.data_in(ME_L3L4_L2D4PHI3X2_CM_L3L4_L2D4PHI3X2),
.enable(ME_L3L4_L2D4PHI3X2_CM_L3L4_L2D4PHI3X2_wr_en),
.number_out(CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4),
.start(ME_L3L4_L2D4PHI3X2_start),
.done(CM_L3L4_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D4PHI4X1_CM_L3L4_L2D4PHI4X1;
wire ME_L3L4_L2D4PHI4X1_CM_L3L4_L2D4PHI4X1_wr_en;
wire [5:0] CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI4X1(
.data_in(ME_L3L4_L2D4PHI4X1_CM_L3L4_L2D4PHI4X1),
.enable(ME_L3L4_L2D4PHI4X1_CM_L3L4_L2D4PHI4X1_wr_en),
.number_out(CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4),
.start(ME_L3L4_L2D4PHI4X1_start),
.done(CM_L3L4_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L2D4PHI4X2_CM_L3L4_L2D4PHI4X2;
wire ME_L3L4_L2D4PHI4X2_CM_L3L4_L2D4PHI4X2_wr_en;
wire [5:0] CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4_number;
wire [8:0] CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4_read_add;
wire [11:0] CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4;
CandidateMatch  CM_L3L4_L2D4PHI4X2(
.data_in(ME_L3L4_L2D4PHI4X2_CM_L3L4_L2D4PHI4X2),
.enable(ME_L3L4_L2D4PHI4X2_CM_L3L4_L2D4PHI4X2_wr_en),
.number_out(CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4_number),
.read_add(CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4_read_add),
.data_out(CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4),
.start(ME_L3L4_L2D4PHI4X2_start),
.done(CM_L3L4_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L2D4_L3L4_AP_L3L4_L2D4;
wire PR_L2D4_L3L4_AP_L3L4_L2D4_wr_en;
wire [8:0] AP_L3L4_L2D4_MC_L3L4_L2D4_read_add;
wire [55:0] AP_L3L4_L2D4_MC_L3L4_L2D4;
AllProj  AP_L3L4_L2D4(
.data_in(PR_L2D4_L3L4_AP_L3L4_L2D4),
.enable(PR_L2D4_L3L4_AP_L3L4_L2D4_wr_en),
.read_add(AP_L3L4_L2D4_MC_L3L4_L2D4_read_add),
.data_out(AP_L3L4_L2D4_MC_L3L4_L2D4),
.start(PR_L2D4_L3L4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L2D4_AS_L2D4n3;
wire VMR_L2D4_AS_L2D4n3_wr_en;
wire [10:0] AS_L2D4n3_MC_L3L4_L2D4_read_add;
wire [35:0] AS_L2D4n3_MC_L3L4_L2D4;
AllStubs  AS_L2D4n3(
.data_in(VMR_L2D4_AS_L2D4n3),
.enable(VMR_L2D4_AS_L2D4n3_wr_en),
.read_add_MC(AS_L2D4n3_MC_L3L4_L2D4_read_add),
.data_out_MC(AS_L2D4n3_MC_L3L4_L2D4),
.start(VMR_L2D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D3PHI1X1_CM_L3L4_L5D3PHI1X1;
wire ME_L3L4_L5D3PHI1X1_CM_L3L4_L5D3PHI1X1_wr_en;
wire [5:0] CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI1X1(
.data_in(ME_L3L4_L5D3PHI1X1_CM_L3L4_L5D3PHI1X1),
.enable(ME_L3L4_L5D3PHI1X1_CM_L3L4_L5D3PHI1X1_wr_en),
.number_out(CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3),
.start(ME_L3L4_L5D3PHI1X1_start),
.done(CM_L3L4_L5D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D3PHI1X2_CM_L3L4_L5D3PHI1X2;
wire ME_L3L4_L5D3PHI1X2_CM_L3L4_L5D3PHI1X2_wr_en;
wire [5:0] CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI1X2(
.data_in(ME_L3L4_L5D3PHI1X2_CM_L3L4_L5D3PHI1X2),
.enable(ME_L3L4_L5D3PHI1X2_CM_L3L4_L5D3PHI1X2_wr_en),
.number_out(CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3),
.start(ME_L3L4_L5D3PHI1X2_start),
.done(CM_L3L4_L5D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D3PHI2X1_CM_L3L4_L5D3PHI2X1;
wire ME_L3L4_L5D3PHI2X1_CM_L3L4_L5D3PHI2X1_wr_en;
wire [5:0] CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI2X1(
.data_in(ME_L3L4_L5D3PHI2X1_CM_L3L4_L5D3PHI2X1),
.enable(ME_L3L4_L5D3PHI2X1_CM_L3L4_L5D3PHI2X1_wr_en),
.number_out(CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3),
.start(ME_L3L4_L5D3PHI2X1_start),
.done(CM_L3L4_L5D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D3PHI2X2_CM_L3L4_L5D3PHI2X2;
wire ME_L3L4_L5D3PHI2X2_CM_L3L4_L5D3PHI2X2_wr_en;
wire [5:0] CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI2X2(
.data_in(ME_L3L4_L5D3PHI2X2_CM_L3L4_L5D3PHI2X2),
.enable(ME_L3L4_L5D3PHI2X2_CM_L3L4_L5D3PHI2X2_wr_en),
.number_out(CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3),
.start(ME_L3L4_L5D3PHI2X2_start),
.done(CM_L3L4_L5D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D3PHI3X1_CM_L3L4_L5D3PHI3X1;
wire ME_L3L4_L5D3PHI3X1_CM_L3L4_L5D3PHI3X1_wr_en;
wire [5:0] CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI3X1(
.data_in(ME_L3L4_L5D3PHI3X1_CM_L3L4_L5D3PHI3X1),
.enable(ME_L3L4_L5D3PHI3X1_CM_L3L4_L5D3PHI3X1_wr_en),
.number_out(CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3),
.start(ME_L3L4_L5D3PHI3X1_start),
.done(CM_L3L4_L5D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D3PHI3X2_CM_L3L4_L5D3PHI3X2;
wire ME_L3L4_L5D3PHI3X2_CM_L3L4_L5D3PHI3X2_wr_en;
wire [5:0] CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3_number;
wire [8:0] CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3_read_add;
wire [11:0] CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3;
CandidateMatch  CM_L3L4_L5D3PHI3X2(
.data_in(ME_L3L4_L5D3PHI3X2_CM_L3L4_L5D3PHI3X2),
.enable(ME_L3L4_L5D3PHI3X2_CM_L3L4_L5D3PHI3X2_wr_en),
.number_out(CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3_number),
.read_add(CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3_read_add),
.data_out(CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3),
.start(ME_L3L4_L5D3PHI3X2_start),
.done(CM_L3L4_L5D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L5D3_L3L4_AP_L3L4_L5D3;
wire PR_L5D3_L3L4_AP_L3L4_L5D3_wr_en;
wire [8:0] AP_L3L4_L5D3_MC_L3L4_L5D3_read_add;
wire [55:0] AP_L3L4_L5D3_MC_L3L4_L5D3;
AllProj #(1'b0,1'b0) AP_L3L4_L5D3(
.data_in(PR_L5D3_L3L4_AP_L3L4_L5D3),
.enable(PR_L5D3_L3L4_AP_L3L4_L5D3_wr_en),
.read_add(AP_L3L4_L5D3_MC_L3L4_L5D3_read_add),
.data_out(AP_L3L4_L5D3_MC_L3L4_L5D3),
.start(PR_L5D3_L3L4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L5D3_AS_L5D3n3;
wire VMR_L5D3_AS_L5D3n3_wr_en;
wire [10:0] AS_L5D3n3_MC_L3L4_L5D3_read_add;
wire [35:0] AS_L5D3n3_MC_L3L4_L5D3;
AllStubs  AS_L5D3n3(
.data_in(VMR_L5D3_AS_L5D3n3),
.enable(VMR_L5D3_AS_L5D3n3_wr_en),
.read_add_MC(AS_L5D3n3_MC_L3L4_L5D3_read_add),
.data_out_MC(AS_L5D3n3_MC_L3L4_L5D3),
.start(VMR_L5D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D4PHI1X1_CM_L3L4_L5D4PHI1X1;
wire ME_L3L4_L5D4PHI1X1_CM_L3L4_L5D4PHI1X1_wr_en;
wire [5:0] CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI1X1(
.data_in(ME_L3L4_L5D4PHI1X1_CM_L3L4_L5D4PHI1X1),
.enable(ME_L3L4_L5D4PHI1X1_CM_L3L4_L5D4PHI1X1_wr_en),
.number_out(CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4),
.start(ME_L3L4_L5D4PHI1X1_start),
.done(CM_L3L4_L5D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D4PHI1X2_CM_L3L4_L5D4PHI1X2;
wire ME_L3L4_L5D4PHI1X2_CM_L3L4_L5D4PHI1X2_wr_en;
wire [5:0] CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI1X2(
.data_in(ME_L3L4_L5D4PHI1X2_CM_L3L4_L5D4PHI1X2),
.enable(ME_L3L4_L5D4PHI1X2_CM_L3L4_L5D4PHI1X2_wr_en),
.number_out(CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4),
.start(ME_L3L4_L5D4PHI1X2_start),
.done(CM_L3L4_L5D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D4PHI2X1_CM_L3L4_L5D4PHI2X1;
wire ME_L3L4_L5D4PHI2X1_CM_L3L4_L5D4PHI2X1_wr_en;
wire [5:0] CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI2X1(
.data_in(ME_L3L4_L5D4PHI2X1_CM_L3L4_L5D4PHI2X1),
.enable(ME_L3L4_L5D4PHI2X1_CM_L3L4_L5D4PHI2X1_wr_en),
.number_out(CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4),
.start(ME_L3L4_L5D4PHI2X1_start),
.done(CM_L3L4_L5D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D4PHI2X2_CM_L3L4_L5D4PHI2X2;
wire ME_L3L4_L5D4PHI2X2_CM_L3L4_L5D4PHI2X2_wr_en;
wire [5:0] CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI2X2(
.data_in(ME_L3L4_L5D4PHI2X2_CM_L3L4_L5D4PHI2X2),
.enable(ME_L3L4_L5D4PHI2X2_CM_L3L4_L5D4PHI2X2_wr_en),
.number_out(CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4),
.start(ME_L3L4_L5D4PHI2X2_start),
.done(CM_L3L4_L5D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D4PHI3X1_CM_L3L4_L5D4PHI3X1;
wire ME_L3L4_L5D4PHI3X1_CM_L3L4_L5D4PHI3X1_wr_en;
wire [5:0] CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI3X1(
.data_in(ME_L3L4_L5D4PHI3X1_CM_L3L4_L5D4PHI3X1),
.enable(ME_L3L4_L5D4PHI3X1_CM_L3L4_L5D4PHI3X1_wr_en),
.number_out(CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4),
.start(ME_L3L4_L5D4PHI3X1_start),
.done(CM_L3L4_L5D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L5D4PHI3X2_CM_L3L4_L5D4PHI3X2;
wire ME_L3L4_L5D4PHI3X2_CM_L3L4_L5D4PHI3X2_wr_en;
wire [5:0] CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4_number;
wire [8:0] CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4_read_add;
wire [11:0] CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4;
CandidateMatch  CM_L3L4_L5D4PHI3X2(
.data_in(ME_L3L4_L5D4PHI3X2_CM_L3L4_L5D4PHI3X2),
.enable(ME_L3L4_L5D4PHI3X2_CM_L3L4_L5D4PHI3X2_wr_en),
.number_out(CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4_number),
.read_add(CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4_read_add),
.data_out(CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4),
.start(ME_L3L4_L5D4PHI3X2_start),
.done(CM_L3L4_L5D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L5D4_L3L4_AP_L3L4_L5D4;
wire PR_L5D4_L3L4_AP_L3L4_L5D4_wr_en;
wire [8:0] AP_L3L4_L5D4_MC_L3L4_L5D4_read_add;
wire [55:0] AP_L3L4_L5D4_MC_L3L4_L5D4;
AllProj #(1'b0,1'b0) AP_L3L4_L5D4(
.data_in(PR_L5D4_L3L4_AP_L3L4_L5D4),
.enable(PR_L5D4_L3L4_AP_L3L4_L5D4_wr_en),
.read_add(AP_L3L4_L5D4_MC_L3L4_L5D4_read_add),
.data_out(AP_L3L4_L5D4_MC_L3L4_L5D4),
.start(PR_L5D4_L3L4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L5D4_AS_L5D4n2;
wire VMR_L5D4_AS_L5D4n2_wr_en;
wire [10:0] AS_L5D4n2_MC_L3L4_L5D4_read_add;
wire [35:0] AS_L5D4n2_MC_L3L4_L5D4;
AllStubs  AS_L5D4n2(
.data_in(VMR_L5D4_AS_L5D4n2),
.enable(VMR_L5D4_AS_L5D4n2_wr_en),
.read_add_MC(AS_L5D4n2_MC_L3L4_L5D4_read_add),
.data_out_MC(AS_L5D4n2_MC_L3L4_L5D4),
.start(VMR_L5D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D3PHI1X1_CM_L3L4_L6D3PHI1X1;
wire ME_L3L4_L6D3PHI1X1_CM_L3L4_L6D3PHI1X1_wr_en;
wire [5:0] CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI1X1(
.data_in(ME_L3L4_L6D3PHI1X1_CM_L3L4_L6D3PHI1X1),
.enable(ME_L3L4_L6D3PHI1X1_CM_L3L4_L6D3PHI1X1_wr_en),
.number_out(CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3),
.start(ME_L3L4_L6D3PHI1X1_start),
.done(CM_L3L4_L6D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D3PHI1X2_CM_L3L4_L6D3PHI1X2;
wire ME_L3L4_L6D3PHI1X2_CM_L3L4_L6D3PHI1X2_wr_en;
wire [5:0] CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI1X2(
.data_in(ME_L3L4_L6D3PHI1X2_CM_L3L4_L6D3PHI1X2),
.enable(ME_L3L4_L6D3PHI1X2_CM_L3L4_L6D3PHI1X2_wr_en),
.number_out(CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3),
.start(ME_L3L4_L6D3PHI1X2_start),
.done(CM_L3L4_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D3PHI2X1_CM_L3L4_L6D3PHI2X1;
wire ME_L3L4_L6D3PHI2X1_CM_L3L4_L6D3PHI2X1_wr_en;
wire [5:0] CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI2X1(
.data_in(ME_L3L4_L6D3PHI2X1_CM_L3L4_L6D3PHI2X1),
.enable(ME_L3L4_L6D3PHI2X1_CM_L3L4_L6D3PHI2X1_wr_en),
.number_out(CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3),
.start(ME_L3L4_L6D3PHI2X1_start),
.done(CM_L3L4_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D3PHI2X2_CM_L3L4_L6D3PHI2X2;
wire ME_L3L4_L6D3PHI2X2_CM_L3L4_L6D3PHI2X2_wr_en;
wire [5:0] CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI2X2(
.data_in(ME_L3L4_L6D3PHI2X2_CM_L3L4_L6D3PHI2X2),
.enable(ME_L3L4_L6D3PHI2X2_CM_L3L4_L6D3PHI2X2_wr_en),
.number_out(CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3),
.start(ME_L3L4_L6D3PHI2X2_start),
.done(CM_L3L4_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D3PHI3X1_CM_L3L4_L6D3PHI3X1;
wire ME_L3L4_L6D3PHI3X1_CM_L3L4_L6D3PHI3X1_wr_en;
wire [5:0] CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI3X1(
.data_in(ME_L3L4_L6D3PHI3X1_CM_L3L4_L6D3PHI3X1),
.enable(ME_L3L4_L6D3PHI3X1_CM_L3L4_L6D3PHI3X1_wr_en),
.number_out(CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3),
.start(ME_L3L4_L6D3PHI3X1_start),
.done(CM_L3L4_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D3PHI3X2_CM_L3L4_L6D3PHI3X2;
wire ME_L3L4_L6D3PHI3X2_CM_L3L4_L6D3PHI3X2_wr_en;
wire [5:0] CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI3X2(
.data_in(ME_L3L4_L6D3PHI3X2_CM_L3L4_L6D3PHI3X2),
.enable(ME_L3L4_L6D3PHI3X2_CM_L3L4_L6D3PHI3X2_wr_en),
.number_out(CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3),
.start(ME_L3L4_L6D3PHI3X2_start),
.done(CM_L3L4_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D3PHI4X1_CM_L3L4_L6D3PHI4X1;
wire ME_L3L4_L6D3PHI4X1_CM_L3L4_L6D3PHI4X1_wr_en;
wire [5:0] CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI4X1(
.data_in(ME_L3L4_L6D3PHI4X1_CM_L3L4_L6D3PHI4X1),
.enable(ME_L3L4_L6D3PHI4X1_CM_L3L4_L6D3PHI4X1_wr_en),
.number_out(CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3),
.start(ME_L3L4_L6D3PHI4X1_start),
.done(CM_L3L4_L6D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D3PHI4X2_CM_L3L4_L6D3PHI4X2;
wire ME_L3L4_L6D3PHI4X2_CM_L3L4_L6D3PHI4X2_wr_en;
wire [5:0] CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3_number;
wire [8:0] CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3_read_add;
wire [11:0] CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3;
CandidateMatch  CM_L3L4_L6D3PHI4X2(
.data_in(ME_L3L4_L6D3PHI4X2_CM_L3L4_L6D3PHI4X2),
.enable(ME_L3L4_L6D3PHI4X2_CM_L3L4_L6D3PHI4X2_wr_en),
.number_out(CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3_number),
.read_add(CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3_read_add),
.data_out(CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3),
.start(ME_L3L4_L6D3PHI4X2_start),
.done(CM_L3L4_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L6D3_L3L4_AP_L3L4_L6D3;
wire PR_L6D3_L3L4_AP_L3L4_L6D3_wr_en;
wire [8:0] AP_L3L4_L6D3_MC_L3L4_L6D3_read_add;
wire [55:0] AP_L3L4_L6D3_MC_L3L4_L6D3;
AllProj #(1'b0,1'b0) AP_L3L4_L6D3(
.data_in(PR_L6D3_L3L4_AP_L3L4_L6D3),
.enable(PR_L6D3_L3L4_AP_L3L4_L6D3_wr_en),
.read_add(AP_L3L4_L6D3_MC_L3L4_L6D3_read_add),
.data_out(AP_L3L4_L6D3_MC_L3L4_L6D3),
.start(PR_L6D3_L3L4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L6D3_AS_L6D3n2;
wire VMR_L6D3_AS_L6D3n2_wr_en;
wire [10:0] AS_L6D3n2_MC_L3L4_L6D3_read_add;
wire [35:0] AS_L6D3n2_MC_L3L4_L6D3;
AllStubs  AS_L6D3n2(
.data_in(VMR_L6D3_AS_L6D3n2),
.enable(VMR_L6D3_AS_L6D3n2_wr_en),
.read_add_MC(AS_L6D3n2_MC_L3L4_L6D3_read_add),
.data_out_MC(AS_L6D3n2_MC_L3L4_L6D3),
.start(VMR_L6D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D4PHI1X1_CM_L3L4_L6D4PHI1X1;
wire ME_L3L4_L6D4PHI1X1_CM_L3L4_L6D4PHI1X1_wr_en;
wire [5:0] CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI1X1(
.data_in(ME_L3L4_L6D4PHI1X1_CM_L3L4_L6D4PHI1X1),
.enable(ME_L3L4_L6D4PHI1X1_CM_L3L4_L6D4PHI1X1_wr_en),
.number_out(CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4),
.start(ME_L3L4_L6D4PHI1X1_start),
.done(CM_L3L4_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D4PHI1X2_CM_L3L4_L6D4PHI1X2;
wire ME_L3L4_L6D4PHI1X2_CM_L3L4_L6D4PHI1X2_wr_en;
wire [5:0] CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI1X2(
.data_in(ME_L3L4_L6D4PHI1X2_CM_L3L4_L6D4PHI1X2),
.enable(ME_L3L4_L6D4PHI1X2_CM_L3L4_L6D4PHI1X2_wr_en),
.number_out(CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4),
.start(ME_L3L4_L6D4PHI1X2_start),
.done(CM_L3L4_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D4PHI2X1_CM_L3L4_L6D4PHI2X1;
wire ME_L3L4_L6D4PHI2X1_CM_L3L4_L6D4PHI2X1_wr_en;
wire [5:0] CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI2X1(
.data_in(ME_L3L4_L6D4PHI2X1_CM_L3L4_L6D4PHI2X1),
.enable(ME_L3L4_L6D4PHI2X1_CM_L3L4_L6D4PHI2X1_wr_en),
.number_out(CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4),
.start(ME_L3L4_L6D4PHI2X1_start),
.done(CM_L3L4_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D4PHI2X2_CM_L3L4_L6D4PHI2X2;
wire ME_L3L4_L6D4PHI2X2_CM_L3L4_L6D4PHI2X2_wr_en;
wire [5:0] CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI2X2(
.data_in(ME_L3L4_L6D4PHI2X2_CM_L3L4_L6D4PHI2X2),
.enable(ME_L3L4_L6D4PHI2X2_CM_L3L4_L6D4PHI2X2_wr_en),
.number_out(CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4),
.start(ME_L3L4_L6D4PHI2X2_start),
.done(CM_L3L4_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D4PHI3X1_CM_L3L4_L6D4PHI3X1;
wire ME_L3L4_L6D4PHI3X1_CM_L3L4_L6D4PHI3X1_wr_en;
wire [5:0] CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI3X1(
.data_in(ME_L3L4_L6D4PHI3X1_CM_L3L4_L6D4PHI3X1),
.enable(ME_L3L4_L6D4PHI3X1_CM_L3L4_L6D4PHI3X1_wr_en),
.number_out(CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4),
.start(ME_L3L4_L6D4PHI3X1_start),
.done(CM_L3L4_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D4PHI3X2_CM_L3L4_L6D4PHI3X2;
wire ME_L3L4_L6D4PHI3X2_CM_L3L4_L6D4PHI3X2_wr_en;
wire [5:0] CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI3X2(
.data_in(ME_L3L4_L6D4PHI3X2_CM_L3L4_L6D4PHI3X2),
.enable(ME_L3L4_L6D4PHI3X2_CM_L3L4_L6D4PHI3X2_wr_en),
.number_out(CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4),
.start(ME_L3L4_L6D4PHI3X2_start),
.done(CM_L3L4_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D4PHI4X1_CM_L3L4_L6D4PHI4X1;
wire ME_L3L4_L6D4PHI4X1_CM_L3L4_L6D4PHI4X1_wr_en;
wire [5:0] CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI4X1(
.data_in(ME_L3L4_L6D4PHI4X1_CM_L3L4_L6D4PHI4X1),
.enable(ME_L3L4_L6D4PHI4X1_CM_L3L4_L6D4PHI4X1_wr_en),
.number_out(CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4),
.start(ME_L3L4_L6D4PHI4X1_start),
.done(CM_L3L4_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L3L4_L6D4PHI4X2_CM_L3L4_L6D4PHI4X2;
wire ME_L3L4_L6D4PHI4X2_CM_L3L4_L6D4PHI4X2_wr_en;
wire [5:0] CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4_number;
wire [8:0] CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4_read_add;
wire [11:0] CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4;
CandidateMatch  CM_L3L4_L6D4PHI4X2(
.data_in(ME_L3L4_L6D4PHI4X2_CM_L3L4_L6D4PHI4X2),
.enable(ME_L3L4_L6D4PHI4X2_CM_L3L4_L6D4PHI4X2_wr_en),
.number_out(CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4_number),
.read_add(CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4_read_add),
.data_out(CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4),
.start(ME_L3L4_L6D4PHI4X2_start),
.done(CM_L3L4_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L6D4_L3L4_AP_L3L4_L6D4;
wire PR_L6D4_L3L4_AP_L3L4_L6D4_wr_en;
wire [8:0] AP_L3L4_L6D4_MC_L3L4_L6D4_read_add;
wire [55:0] AP_L3L4_L6D4_MC_L3L4_L6D4;
AllProj #(1'b0,1'b0) AP_L3L4_L6D4(
.data_in(PR_L6D4_L3L4_AP_L3L4_L6D4),
.enable(PR_L6D4_L3L4_AP_L3L4_L6D4_wr_en),
.read_add(AP_L3L4_L6D4_MC_L3L4_L6D4_read_add),
.data_out(AP_L3L4_L6D4_MC_L3L4_L6D4),
.start(PR_L6D4_L3L4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L6D4_AS_L6D4n3;
wire VMR_L6D4_AS_L6D4n3_wr_en;
wire [10:0] AS_L6D4n3_MC_L3L4_L6D4_read_add;
wire [35:0] AS_L6D4n3_MC_L3L4_L6D4;
AllStubs  AS_L6D4n3(
.data_in(VMR_L6D4_AS_L6D4n3),
.enable(VMR_L6D4_AS_L6D4n3_wr_en),
.read_add_MC(AS_L6D4n3_MC_L3L4_L6D4_read_add),
.data_out_MC(AS_L6D4n3_MC_L3L4_L6D4),
.start(VMR_L6D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D3PHI1X1_CM_L5L6_L1D3PHI1X1;
wire ME_L5L6_L1D3PHI1X1_CM_L5L6_L1D3PHI1X1_wr_en;
wire [5:0] CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI1X1(
.data_in(ME_L5L6_L1D3PHI1X1_CM_L5L6_L1D3PHI1X1),
.enable(ME_L5L6_L1D3PHI1X1_CM_L5L6_L1D3PHI1X1_wr_en),
.number_out(CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3),
.start(ME_L5L6_L1D3PHI1X1_start),
.done(CM_L5L6_L1D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D3PHI1X2_CM_L5L6_L1D3PHI1X2;
wire ME_L5L6_L1D3PHI1X2_CM_L5L6_L1D3PHI1X2_wr_en;
wire [5:0] CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI1X2(
.data_in(ME_L5L6_L1D3PHI1X2_CM_L5L6_L1D3PHI1X2),
.enable(ME_L5L6_L1D3PHI1X2_CM_L5L6_L1D3PHI1X2_wr_en),
.number_out(CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3),
.start(ME_L5L6_L1D3PHI1X2_start),
.done(CM_L5L6_L1D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D3PHI2X1_CM_L5L6_L1D3PHI2X1;
wire ME_L5L6_L1D3PHI2X1_CM_L5L6_L1D3PHI2X1_wr_en;
wire [5:0] CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI2X1(
.data_in(ME_L5L6_L1D3PHI2X1_CM_L5L6_L1D3PHI2X1),
.enable(ME_L5L6_L1D3PHI2X1_CM_L5L6_L1D3PHI2X1_wr_en),
.number_out(CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3),
.start(ME_L5L6_L1D3PHI2X1_start),
.done(CM_L5L6_L1D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D3PHI2X2_CM_L5L6_L1D3PHI2X2;
wire ME_L5L6_L1D3PHI2X2_CM_L5L6_L1D3PHI2X2_wr_en;
wire [5:0] CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI2X2(
.data_in(ME_L5L6_L1D3PHI2X2_CM_L5L6_L1D3PHI2X2),
.enable(ME_L5L6_L1D3PHI2X2_CM_L5L6_L1D3PHI2X2_wr_en),
.number_out(CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3),
.start(ME_L5L6_L1D3PHI2X2_start),
.done(CM_L5L6_L1D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D3PHI3X1_CM_L5L6_L1D3PHI3X1;
wire ME_L5L6_L1D3PHI3X1_CM_L5L6_L1D3PHI3X1_wr_en;
wire [5:0] CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI3X1(
.data_in(ME_L5L6_L1D3PHI3X1_CM_L5L6_L1D3PHI3X1),
.enable(ME_L5L6_L1D3PHI3X1_CM_L5L6_L1D3PHI3X1_wr_en),
.number_out(CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3),
.start(ME_L5L6_L1D3PHI3X1_start),
.done(CM_L5L6_L1D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D3PHI3X2_CM_L5L6_L1D3PHI3X2;
wire ME_L5L6_L1D3PHI3X2_CM_L5L6_L1D3PHI3X2_wr_en;
wire [5:0] CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3_number;
wire [8:0] CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3_read_add;
wire [11:0] CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3;
CandidateMatch  CM_L5L6_L1D3PHI3X2(
.data_in(ME_L5L6_L1D3PHI3X2_CM_L5L6_L1D3PHI3X2),
.enable(ME_L5L6_L1D3PHI3X2_CM_L5L6_L1D3PHI3X2_wr_en),
.number_out(CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3_number),
.read_add(CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3_read_add),
.data_out(CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3),
.start(ME_L5L6_L1D3PHI3X2_start),
.done(CM_L5L6_L1D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L1D3_L5L6_AP_L5L6_L1D3;
wire PR_L1D3_L5L6_AP_L5L6_L1D3_wr_en;
wire [8:0] AP_L5L6_L1D3_MC_L5L6_L1D3_read_add;
wire [55:0] AP_L5L6_L1D3_MC_L5L6_L1D3;
AllProj  AP_L5L6_L1D3(
.data_in(PR_L1D3_L5L6_AP_L5L6_L1D3),
.enable(PR_L1D3_L5L6_AP_L5L6_L1D3_wr_en),
.read_add(AP_L5L6_L1D3_MC_L5L6_L1D3_read_add),
.data_out(AP_L5L6_L1D3_MC_L5L6_L1D3),
.start(PR_L1D3_L5L6_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L1D3_AS_L1D3n4;
wire VMR_L1D3_AS_L1D3n4_wr_en;
wire [10:0] AS_L1D3n4_MC_L5L6_L1D3_read_add;
wire [35:0] AS_L1D3n4_MC_L5L6_L1D3;
AllStubs  AS_L1D3n4(
.data_in(VMR_L1D3_AS_L1D3n4),
.enable(VMR_L1D3_AS_L1D3n4_wr_en),
.read_add_MC(AS_L1D3n4_MC_L5L6_L1D3_read_add),
.data_out_MC(AS_L1D3n4_MC_L5L6_L1D3),
.start(VMR_L1D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D4PHI1X1_CM_L5L6_L1D4PHI1X1;
wire ME_L5L6_L1D4PHI1X1_CM_L5L6_L1D4PHI1X1_wr_en;
wire [5:0] CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI1X1(
.data_in(ME_L5L6_L1D4PHI1X1_CM_L5L6_L1D4PHI1X1),
.enable(ME_L5L6_L1D4PHI1X1_CM_L5L6_L1D4PHI1X1_wr_en),
.number_out(CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4),
.start(ME_L5L6_L1D4PHI1X1_start),
.done(CM_L5L6_L1D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D4PHI1X2_CM_L5L6_L1D4PHI1X2;
wire ME_L5L6_L1D4PHI1X2_CM_L5L6_L1D4PHI1X2_wr_en;
wire [5:0] CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI1X2(
.data_in(ME_L5L6_L1D4PHI1X2_CM_L5L6_L1D4PHI1X2),
.enable(ME_L5L6_L1D4PHI1X2_CM_L5L6_L1D4PHI1X2_wr_en),
.number_out(CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4),
.start(ME_L5L6_L1D4PHI1X2_start),
.done(CM_L5L6_L1D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D4PHI2X1_CM_L5L6_L1D4PHI2X1;
wire ME_L5L6_L1D4PHI2X1_CM_L5L6_L1D4PHI2X1_wr_en;
wire [5:0] CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI2X1(
.data_in(ME_L5L6_L1D4PHI2X1_CM_L5L6_L1D4PHI2X1),
.enable(ME_L5L6_L1D4PHI2X1_CM_L5L6_L1D4PHI2X1_wr_en),
.number_out(CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4),
.start(ME_L5L6_L1D4PHI2X1_start),
.done(CM_L5L6_L1D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D4PHI2X2_CM_L5L6_L1D4PHI2X2;
wire ME_L5L6_L1D4PHI2X2_CM_L5L6_L1D4PHI2X2_wr_en;
wire [5:0] CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI2X2(
.data_in(ME_L5L6_L1D4PHI2X2_CM_L5L6_L1D4PHI2X2),
.enable(ME_L5L6_L1D4PHI2X2_CM_L5L6_L1D4PHI2X2_wr_en),
.number_out(CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4),
.start(ME_L5L6_L1D4PHI2X2_start),
.done(CM_L5L6_L1D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D4PHI3X1_CM_L5L6_L1D4PHI3X1;
wire ME_L5L6_L1D4PHI3X1_CM_L5L6_L1D4PHI3X1_wr_en;
wire [5:0] CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI3X1(
.data_in(ME_L5L6_L1D4PHI3X1_CM_L5L6_L1D4PHI3X1),
.enable(ME_L5L6_L1D4PHI3X1_CM_L5L6_L1D4PHI3X1_wr_en),
.number_out(CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4),
.start(ME_L5L6_L1D4PHI3X1_start),
.done(CM_L5L6_L1D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L1D4PHI3X2_CM_L5L6_L1D4PHI3X2;
wire ME_L5L6_L1D4PHI3X2_CM_L5L6_L1D4PHI3X2_wr_en;
wire [5:0] CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4_number;
wire [8:0] CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4_read_add;
wire [11:0] CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4;
CandidateMatch  CM_L5L6_L1D4PHI3X2(
.data_in(ME_L5L6_L1D4PHI3X2_CM_L5L6_L1D4PHI3X2),
.enable(ME_L5L6_L1D4PHI3X2_CM_L5L6_L1D4PHI3X2_wr_en),
.number_out(CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4_number),
.read_add(CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4_read_add),
.data_out(CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4),
.start(ME_L5L6_L1D4PHI3X2_start),
.done(CM_L5L6_L1D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L1D4_L5L6_AP_L5L6_L1D4;
wire PR_L1D4_L5L6_AP_L5L6_L1D4_wr_en;
wire [8:0] AP_L5L6_L1D4_MC_L5L6_L1D4_read_add;
wire [55:0] AP_L5L6_L1D4_MC_L5L6_L1D4;
AllProj  AP_L5L6_L1D4(
.data_in(PR_L1D4_L5L6_AP_L5L6_L1D4),
.enable(PR_L1D4_L5L6_AP_L5L6_L1D4_wr_en),
.read_add(AP_L5L6_L1D4_MC_L5L6_L1D4_read_add),
.data_out(AP_L5L6_L1D4_MC_L5L6_L1D4),
.start(PR_L1D4_L5L6_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L1D4_AS_L1D4n3;
wire VMR_L1D4_AS_L1D4n3_wr_en;
wire [10:0] AS_L1D4n3_MC_L5L6_L1D4_read_add;
wire [35:0] AS_L1D4n3_MC_L5L6_L1D4;
AllStubs  AS_L1D4n3(
.data_in(VMR_L1D4_AS_L1D4n3),
.enable(VMR_L1D4_AS_L1D4n3_wr_en),
.read_add_MC(AS_L1D4n3_MC_L5L6_L1D4_read_add),
.data_out_MC(AS_L1D4n3_MC_L5L6_L1D4),
.start(VMR_L1D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D3PHI1X1_CM_L5L6_L2D3PHI1X1;
wire ME_L5L6_L2D3PHI1X1_CM_L5L6_L2D3PHI1X1_wr_en;
wire [5:0] CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI1X1(
.data_in(ME_L5L6_L2D3PHI1X1_CM_L5L6_L2D3PHI1X1),
.enable(ME_L5L6_L2D3PHI1X1_CM_L5L6_L2D3PHI1X1_wr_en),
.number_out(CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3),
.start(ME_L5L6_L2D3PHI1X1_start),
.done(CM_L5L6_L2D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D3PHI1X2_CM_L5L6_L2D3PHI1X2;
wire ME_L5L6_L2D3PHI1X2_CM_L5L6_L2D3PHI1X2_wr_en;
wire [5:0] CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI1X2(
.data_in(ME_L5L6_L2D3PHI1X2_CM_L5L6_L2D3PHI1X2),
.enable(ME_L5L6_L2D3PHI1X2_CM_L5L6_L2D3PHI1X2_wr_en),
.number_out(CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3),
.start(ME_L5L6_L2D3PHI1X2_start),
.done(CM_L5L6_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D3PHI2X1_CM_L5L6_L2D3PHI2X1;
wire ME_L5L6_L2D3PHI2X1_CM_L5L6_L2D3PHI2X1_wr_en;
wire [5:0] CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI2X1(
.data_in(ME_L5L6_L2D3PHI2X1_CM_L5L6_L2D3PHI2X1),
.enable(ME_L5L6_L2D3PHI2X1_CM_L5L6_L2D3PHI2X1_wr_en),
.number_out(CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3),
.start(ME_L5L6_L2D3PHI2X1_start),
.done(CM_L5L6_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D3PHI2X2_CM_L5L6_L2D3PHI2X2;
wire ME_L5L6_L2D3PHI2X2_CM_L5L6_L2D3PHI2X2_wr_en;
wire [5:0] CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI2X2(
.data_in(ME_L5L6_L2D3PHI2X2_CM_L5L6_L2D3PHI2X2),
.enable(ME_L5L6_L2D3PHI2X2_CM_L5L6_L2D3PHI2X2_wr_en),
.number_out(CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3),
.start(ME_L5L6_L2D3PHI2X2_start),
.done(CM_L5L6_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D3PHI3X1_CM_L5L6_L2D3PHI3X1;
wire ME_L5L6_L2D3PHI3X1_CM_L5L6_L2D3PHI3X1_wr_en;
wire [5:0] CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI3X1(
.data_in(ME_L5L6_L2D3PHI3X1_CM_L5L6_L2D3PHI3X1),
.enable(ME_L5L6_L2D3PHI3X1_CM_L5L6_L2D3PHI3X1_wr_en),
.number_out(CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3),
.start(ME_L5L6_L2D3PHI3X1_start),
.done(CM_L5L6_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D3PHI3X2_CM_L5L6_L2D3PHI3X2;
wire ME_L5L6_L2D3PHI3X2_CM_L5L6_L2D3PHI3X2_wr_en;
wire [5:0] CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI3X2(
.data_in(ME_L5L6_L2D3PHI3X2_CM_L5L6_L2D3PHI3X2),
.enable(ME_L5L6_L2D3PHI3X2_CM_L5L6_L2D3PHI3X2_wr_en),
.number_out(CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3),
.start(ME_L5L6_L2D3PHI3X2_start),
.done(CM_L5L6_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D3PHI4X1_CM_L5L6_L2D3PHI4X1;
wire ME_L5L6_L2D3PHI4X1_CM_L5L6_L2D3PHI4X1_wr_en;
wire [5:0] CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI4X1(
.data_in(ME_L5L6_L2D3PHI4X1_CM_L5L6_L2D3PHI4X1),
.enable(ME_L5L6_L2D3PHI4X1_CM_L5L6_L2D3PHI4X1_wr_en),
.number_out(CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3),
.start(ME_L5L6_L2D3PHI4X1_start),
.done(CM_L5L6_L2D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D3PHI4X2_CM_L5L6_L2D3PHI4X2;
wire ME_L5L6_L2D3PHI4X2_CM_L5L6_L2D3PHI4X2_wr_en;
wire [5:0] CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3_number;
wire [8:0] CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3_read_add;
wire [11:0] CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3;
CandidateMatch  CM_L5L6_L2D3PHI4X2(
.data_in(ME_L5L6_L2D3PHI4X2_CM_L5L6_L2D3PHI4X2),
.enable(ME_L5L6_L2D3PHI4X2_CM_L5L6_L2D3PHI4X2_wr_en),
.number_out(CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3_number),
.read_add(CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3_read_add),
.data_out(CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3),
.start(ME_L5L6_L2D3PHI4X2_start),
.done(CM_L5L6_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L2D3_L5L6_AP_L5L6_L2D3;
wire PR_L2D3_L5L6_AP_L5L6_L2D3_wr_en;
wire [8:0] AP_L5L6_L2D3_MC_L5L6_L2D3_read_add;
wire [55:0] AP_L5L6_L2D3_MC_L5L6_L2D3;
AllProj  AP_L5L6_L2D3(
.data_in(PR_L2D3_L5L6_AP_L5L6_L2D3),
.enable(PR_L2D3_L5L6_AP_L5L6_L2D3_wr_en),
.read_add(AP_L5L6_L2D3_MC_L5L6_L2D3_read_add),
.data_out(AP_L5L6_L2D3_MC_L5L6_L2D3),
.start(PR_L2D3_L5L6_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L2D3_AS_L2D3n3;
wire VMR_L2D3_AS_L2D3n3_wr_en;
wire [10:0] AS_L2D3n3_MC_L5L6_L2D3_read_add;
wire [35:0] AS_L2D3n3_MC_L5L6_L2D3;
AllStubs  AS_L2D3n3(
.data_in(VMR_L2D3_AS_L2D3n3),
.enable(VMR_L2D3_AS_L2D3n3_wr_en),
.read_add_MC(AS_L2D3n3_MC_L5L6_L2D3_read_add),
.data_out_MC(AS_L2D3n3_MC_L5L6_L2D3),
.start(VMR_L2D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D4PHI1X1_CM_L5L6_L2D4PHI1X1;
wire ME_L5L6_L2D4PHI1X1_CM_L5L6_L2D4PHI1X1_wr_en;
wire [5:0] CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI1X1(
.data_in(ME_L5L6_L2D4PHI1X1_CM_L5L6_L2D4PHI1X1),
.enable(ME_L5L6_L2D4PHI1X1_CM_L5L6_L2D4PHI1X1_wr_en),
.number_out(CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4),
.start(ME_L5L6_L2D4PHI1X1_start),
.done(CM_L5L6_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D4PHI1X2_CM_L5L6_L2D4PHI1X2;
wire ME_L5L6_L2D4PHI1X2_CM_L5L6_L2D4PHI1X2_wr_en;
wire [5:0] CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI1X2(
.data_in(ME_L5L6_L2D4PHI1X2_CM_L5L6_L2D4PHI1X2),
.enable(ME_L5L6_L2D4PHI1X2_CM_L5L6_L2D4PHI1X2_wr_en),
.number_out(CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4),
.start(ME_L5L6_L2D4PHI1X2_start),
.done(CM_L5L6_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D4PHI2X1_CM_L5L6_L2D4PHI2X1;
wire ME_L5L6_L2D4PHI2X1_CM_L5L6_L2D4PHI2X1_wr_en;
wire [5:0] CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI2X1(
.data_in(ME_L5L6_L2D4PHI2X1_CM_L5L6_L2D4PHI2X1),
.enable(ME_L5L6_L2D4PHI2X1_CM_L5L6_L2D4PHI2X1_wr_en),
.number_out(CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4),
.start(ME_L5L6_L2D4PHI2X1_start),
.done(CM_L5L6_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D4PHI2X2_CM_L5L6_L2D4PHI2X2;
wire ME_L5L6_L2D4PHI2X2_CM_L5L6_L2D4PHI2X2_wr_en;
wire [5:0] CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI2X2(
.data_in(ME_L5L6_L2D4PHI2X2_CM_L5L6_L2D4PHI2X2),
.enable(ME_L5L6_L2D4PHI2X2_CM_L5L6_L2D4PHI2X2_wr_en),
.number_out(CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4),
.start(ME_L5L6_L2D4PHI2X2_start),
.done(CM_L5L6_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D4PHI3X1_CM_L5L6_L2D4PHI3X1;
wire ME_L5L6_L2D4PHI3X1_CM_L5L6_L2D4PHI3X1_wr_en;
wire [5:0] CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI3X1(
.data_in(ME_L5L6_L2D4PHI3X1_CM_L5L6_L2D4PHI3X1),
.enable(ME_L5L6_L2D4PHI3X1_CM_L5L6_L2D4PHI3X1_wr_en),
.number_out(CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4),
.start(ME_L5L6_L2D4PHI3X1_start),
.done(CM_L5L6_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D4PHI3X2_CM_L5L6_L2D4PHI3X2;
wire ME_L5L6_L2D4PHI3X2_CM_L5L6_L2D4PHI3X2_wr_en;
wire [5:0] CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI3X2(
.data_in(ME_L5L6_L2D4PHI3X2_CM_L5L6_L2D4PHI3X2),
.enable(ME_L5L6_L2D4PHI3X2_CM_L5L6_L2D4PHI3X2_wr_en),
.number_out(CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4),
.start(ME_L5L6_L2D4PHI3X2_start),
.done(CM_L5L6_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D4PHI4X1_CM_L5L6_L2D4PHI4X1;
wire ME_L5L6_L2D4PHI4X1_CM_L5L6_L2D4PHI4X1_wr_en;
wire [5:0] CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI4X1(
.data_in(ME_L5L6_L2D4PHI4X1_CM_L5L6_L2D4PHI4X1),
.enable(ME_L5L6_L2D4PHI4X1_CM_L5L6_L2D4PHI4X1_wr_en),
.number_out(CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4),
.start(ME_L5L6_L2D4PHI4X1_start),
.done(CM_L5L6_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L2D4PHI4X2_CM_L5L6_L2D4PHI4X2;
wire ME_L5L6_L2D4PHI4X2_CM_L5L6_L2D4PHI4X2_wr_en;
wire [5:0] CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4_number;
wire [8:0] CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4_read_add;
wire [11:0] CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4;
CandidateMatch  CM_L5L6_L2D4PHI4X2(
.data_in(ME_L5L6_L2D4PHI4X2_CM_L5L6_L2D4PHI4X2),
.enable(ME_L5L6_L2D4PHI4X2_CM_L5L6_L2D4PHI4X2_wr_en),
.number_out(CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4_number),
.read_add(CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4_read_add),
.data_out(CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4),
.start(ME_L5L6_L2D4PHI4X2_start),
.done(CM_L5L6_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L2D4_L5L6_AP_L5L6_L2D4;
wire PR_L2D4_L5L6_AP_L5L6_L2D4_wr_en;
wire [8:0] AP_L5L6_L2D4_MC_L5L6_L2D4_read_add;
wire [55:0] AP_L5L6_L2D4_MC_L5L6_L2D4;
AllProj  AP_L5L6_L2D4(
.data_in(PR_L2D4_L5L6_AP_L5L6_L2D4),
.enable(PR_L2D4_L5L6_AP_L5L6_L2D4_wr_en),
.read_add(AP_L5L6_L2D4_MC_L5L6_L2D4_read_add),
.data_out(AP_L5L6_L2D4_MC_L5L6_L2D4),
.start(PR_L2D4_L5L6_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L2D4_AS_L2D4n4;
wire VMR_L2D4_AS_L2D4n4_wr_en;
wire [10:0] AS_L2D4n4_MC_L5L6_L2D4_read_add;
wire [35:0] AS_L2D4n4_MC_L5L6_L2D4;
AllStubs  AS_L2D4n4(
.data_in(VMR_L2D4_AS_L2D4n4),
.enable(VMR_L2D4_AS_L2D4n4_wr_en),
.read_add_MC(AS_L2D4n4_MC_L5L6_L2D4_read_add),
.data_out_MC(AS_L2D4n4_MC_L5L6_L2D4),
.start(VMR_L2D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D3PHI1X1_CM_L5L6_L3D3PHI1X1;
wire ME_L5L6_L3D3PHI1X1_CM_L5L6_L3D3PHI1X1_wr_en;
wire [5:0] CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI1X1(
.data_in(ME_L5L6_L3D3PHI1X1_CM_L5L6_L3D3PHI1X1),
.enable(ME_L5L6_L3D3PHI1X1_CM_L5L6_L3D3PHI1X1_wr_en),
.number_out(CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3),
.start(ME_L5L6_L3D3PHI1X1_start),
.done(CM_L5L6_L3D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D3PHI1X2_CM_L5L6_L3D3PHI1X2;
wire ME_L5L6_L3D3PHI1X2_CM_L5L6_L3D3PHI1X2_wr_en;
wire [5:0] CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI1X2(
.data_in(ME_L5L6_L3D3PHI1X2_CM_L5L6_L3D3PHI1X2),
.enable(ME_L5L6_L3D3PHI1X2_CM_L5L6_L3D3PHI1X2_wr_en),
.number_out(CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3),
.start(ME_L5L6_L3D3PHI1X2_start),
.done(CM_L5L6_L3D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D3PHI2X1_CM_L5L6_L3D3PHI2X1;
wire ME_L5L6_L3D3PHI2X1_CM_L5L6_L3D3PHI2X1_wr_en;
wire [5:0] CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI2X1(
.data_in(ME_L5L6_L3D3PHI2X1_CM_L5L6_L3D3PHI2X1),
.enable(ME_L5L6_L3D3PHI2X1_CM_L5L6_L3D3PHI2X1_wr_en),
.number_out(CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3),
.start(ME_L5L6_L3D3PHI2X1_start),
.done(CM_L5L6_L3D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D3PHI2X2_CM_L5L6_L3D3PHI2X2;
wire ME_L5L6_L3D3PHI2X2_CM_L5L6_L3D3PHI2X2_wr_en;
wire [5:0] CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI2X2(
.data_in(ME_L5L6_L3D3PHI2X2_CM_L5L6_L3D3PHI2X2),
.enable(ME_L5L6_L3D3PHI2X2_CM_L5L6_L3D3PHI2X2_wr_en),
.number_out(CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3),
.start(ME_L5L6_L3D3PHI2X2_start),
.done(CM_L5L6_L3D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D3PHI3X1_CM_L5L6_L3D3PHI3X1;
wire ME_L5L6_L3D3PHI3X1_CM_L5L6_L3D3PHI3X1_wr_en;
wire [5:0] CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI3X1(
.data_in(ME_L5L6_L3D3PHI3X1_CM_L5L6_L3D3PHI3X1),
.enable(ME_L5L6_L3D3PHI3X1_CM_L5L6_L3D3PHI3X1_wr_en),
.number_out(CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3),
.start(ME_L5L6_L3D3PHI3X1_start),
.done(CM_L5L6_L3D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D3PHI3X2_CM_L5L6_L3D3PHI3X2;
wire ME_L5L6_L3D3PHI3X2_CM_L5L6_L3D3PHI3X2_wr_en;
wire [5:0] CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3_number;
wire [8:0] CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3_read_add;
wire [11:0] CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3;
CandidateMatch  CM_L5L6_L3D3PHI3X2(
.data_in(ME_L5L6_L3D3PHI3X2_CM_L5L6_L3D3PHI3X2),
.enable(ME_L5L6_L3D3PHI3X2_CM_L5L6_L3D3PHI3X2_wr_en),
.number_out(CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3_number),
.read_add(CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3_read_add),
.data_out(CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3),
.start(ME_L5L6_L3D3PHI3X2_start),
.done(CM_L5L6_L3D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L3D3_L5L6_AP_L5L6_L3D3;
wire PR_L3D3_L5L6_AP_L5L6_L3D3_wr_en;
wire [8:0] AP_L5L6_L3D3_MC_L5L6_L3D3_read_add;
wire [55:0] AP_L5L6_L3D3_MC_L5L6_L3D3;
AllProj  AP_L5L6_L3D3(
.data_in(PR_L3D3_L5L6_AP_L5L6_L3D3),
.enable(PR_L3D3_L5L6_AP_L5L6_L3D3_wr_en),
.read_add(AP_L5L6_L3D3_MC_L5L6_L3D3_read_add),
.data_out(AP_L5L6_L3D3_MC_L5L6_L3D3),
.start(PR_L3D3_L5L6_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L3D3_AS_L3D3n3;
wire VMR_L3D3_AS_L3D3n3_wr_en;
wire [10:0] AS_L3D3n3_MC_L5L6_L3D3_read_add;
wire [35:0] AS_L3D3n3_MC_L5L6_L3D3;
AllStubs  AS_L3D3n3(
.data_in(VMR_L3D3_AS_L3D3n3),
.enable(VMR_L3D3_AS_L3D3n3_wr_en),
.read_add_MC(AS_L3D3n3_MC_L5L6_L3D3_read_add),
.data_out_MC(AS_L3D3n3_MC_L5L6_L3D3),
.start(VMR_L3D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D4PHI1X1_CM_L5L6_L3D4PHI1X1;
wire ME_L5L6_L3D4PHI1X1_CM_L5L6_L3D4PHI1X1_wr_en;
wire [5:0] CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI1X1(
.data_in(ME_L5L6_L3D4PHI1X1_CM_L5L6_L3D4PHI1X1),
.enable(ME_L5L6_L3D4PHI1X1_CM_L5L6_L3D4PHI1X1_wr_en),
.number_out(CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4),
.start(ME_L5L6_L3D4PHI1X1_start),
.done(CM_L5L6_L3D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D4PHI1X2_CM_L5L6_L3D4PHI1X2;
wire ME_L5L6_L3D4PHI1X2_CM_L5L6_L3D4PHI1X2_wr_en;
wire [5:0] CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI1X2(
.data_in(ME_L5L6_L3D4PHI1X2_CM_L5L6_L3D4PHI1X2),
.enable(ME_L5L6_L3D4PHI1X2_CM_L5L6_L3D4PHI1X2_wr_en),
.number_out(CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4),
.start(ME_L5L6_L3D4PHI1X2_start),
.done(CM_L5L6_L3D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D4PHI2X1_CM_L5L6_L3D4PHI2X1;
wire ME_L5L6_L3D4PHI2X1_CM_L5L6_L3D4PHI2X1_wr_en;
wire [5:0] CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI2X1(
.data_in(ME_L5L6_L3D4PHI2X1_CM_L5L6_L3D4PHI2X1),
.enable(ME_L5L6_L3D4PHI2X1_CM_L5L6_L3D4PHI2X1_wr_en),
.number_out(CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4),
.start(ME_L5L6_L3D4PHI2X1_start),
.done(CM_L5L6_L3D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D4PHI2X2_CM_L5L6_L3D4PHI2X2;
wire ME_L5L6_L3D4PHI2X2_CM_L5L6_L3D4PHI2X2_wr_en;
wire [5:0] CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI2X2(
.data_in(ME_L5L6_L3D4PHI2X2_CM_L5L6_L3D4PHI2X2),
.enable(ME_L5L6_L3D4PHI2X2_CM_L5L6_L3D4PHI2X2_wr_en),
.number_out(CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4),
.start(ME_L5L6_L3D4PHI2X2_start),
.done(CM_L5L6_L3D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D4PHI3X1_CM_L5L6_L3D4PHI3X1;
wire ME_L5L6_L3D4PHI3X1_CM_L5L6_L3D4PHI3X1_wr_en;
wire [5:0] CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI3X1(
.data_in(ME_L5L6_L3D4PHI3X1_CM_L5L6_L3D4PHI3X1),
.enable(ME_L5L6_L3D4PHI3X1_CM_L5L6_L3D4PHI3X1_wr_en),
.number_out(CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4),
.start(ME_L5L6_L3D4PHI3X1_start),
.done(CM_L5L6_L3D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L3D4PHI3X2_CM_L5L6_L3D4PHI3X2;
wire ME_L5L6_L3D4PHI3X2_CM_L5L6_L3D4PHI3X2_wr_en;
wire [5:0] CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4_number;
wire [8:0] CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4_read_add;
wire [11:0] CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4;
CandidateMatch  CM_L5L6_L3D4PHI3X2(
.data_in(ME_L5L6_L3D4PHI3X2_CM_L5L6_L3D4PHI3X2),
.enable(ME_L5L6_L3D4PHI3X2_CM_L5L6_L3D4PHI3X2_wr_en),
.number_out(CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4_number),
.read_add(CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4_read_add),
.data_out(CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4),
.start(ME_L5L6_L3D4PHI3X2_start),
.done(CM_L5L6_L3D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L3D4_L5L6_AP_L5L6_L3D4;
wire PR_L3D4_L5L6_AP_L5L6_L3D4_wr_en;
wire [8:0] AP_L5L6_L3D4_MC_L5L6_L3D4_read_add;
wire [55:0] AP_L5L6_L3D4_MC_L5L6_L3D4;
AllProj  AP_L5L6_L3D4(
.data_in(PR_L3D4_L5L6_AP_L5L6_L3D4),
.enable(PR_L3D4_L5L6_AP_L5L6_L3D4_wr_en),
.read_add(AP_L5L6_L3D4_MC_L5L6_L3D4_read_add),
.data_out(AP_L5L6_L3D4_MC_L5L6_L3D4),
.start(PR_L3D4_L5L6_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L3D4_AS_L3D4n2;
wire VMR_L3D4_AS_L3D4n2_wr_en;
wire [10:0] AS_L3D4n2_MC_L5L6_L3D4_read_add;
wire [35:0] AS_L3D4n2_MC_L5L6_L3D4;
AllStubs  AS_L3D4n2(
.data_in(VMR_L3D4_AS_L3D4n2),
.enable(VMR_L3D4_AS_L3D4n2_wr_en),
.read_add_MC(AS_L3D4n2_MC_L5L6_L3D4_read_add),
.data_out_MC(AS_L3D4n2_MC_L5L6_L3D4),
.start(VMR_L3D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D3PHI1X1_CM_L5L6_L4D3PHI1X1;
wire ME_L5L6_L4D3PHI1X1_CM_L5L6_L4D3PHI1X1_wr_en;
wire [5:0] CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI1X1(
.data_in(ME_L5L6_L4D3PHI1X1_CM_L5L6_L4D3PHI1X1),
.enable(ME_L5L6_L4D3PHI1X1_CM_L5L6_L4D3PHI1X1_wr_en),
.number_out(CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3),
.start(ME_L5L6_L4D3PHI1X1_start),
.done(CM_L5L6_L4D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D3PHI1X2_CM_L5L6_L4D3PHI1X2;
wire ME_L5L6_L4D3PHI1X2_CM_L5L6_L4D3PHI1X2_wr_en;
wire [5:0] CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI1X2(
.data_in(ME_L5L6_L4D3PHI1X2_CM_L5L6_L4D3PHI1X2),
.enable(ME_L5L6_L4D3PHI1X2_CM_L5L6_L4D3PHI1X2_wr_en),
.number_out(CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3),
.start(ME_L5L6_L4D3PHI1X2_start),
.done(CM_L5L6_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D3PHI2X1_CM_L5L6_L4D3PHI2X1;
wire ME_L5L6_L4D3PHI2X1_CM_L5L6_L4D3PHI2X1_wr_en;
wire [5:0] CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI2X1(
.data_in(ME_L5L6_L4D3PHI2X1_CM_L5L6_L4D3PHI2X1),
.enable(ME_L5L6_L4D3PHI2X1_CM_L5L6_L4D3PHI2X1_wr_en),
.number_out(CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3),
.start(ME_L5L6_L4D3PHI2X1_start),
.done(CM_L5L6_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D3PHI2X2_CM_L5L6_L4D3PHI2X2;
wire ME_L5L6_L4D3PHI2X2_CM_L5L6_L4D3PHI2X2_wr_en;
wire [5:0] CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI2X2(
.data_in(ME_L5L6_L4D3PHI2X2_CM_L5L6_L4D3PHI2X2),
.enable(ME_L5L6_L4D3PHI2X2_CM_L5L6_L4D3PHI2X2_wr_en),
.number_out(CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3),
.start(ME_L5L6_L4D3PHI2X2_start),
.done(CM_L5L6_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D3PHI3X1_CM_L5L6_L4D3PHI3X1;
wire ME_L5L6_L4D3PHI3X1_CM_L5L6_L4D3PHI3X1_wr_en;
wire [5:0] CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI3X1(
.data_in(ME_L5L6_L4D3PHI3X1_CM_L5L6_L4D3PHI3X1),
.enable(ME_L5L6_L4D3PHI3X1_CM_L5L6_L4D3PHI3X1_wr_en),
.number_out(CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3),
.start(ME_L5L6_L4D3PHI3X1_start),
.done(CM_L5L6_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D3PHI3X2_CM_L5L6_L4D3PHI3X2;
wire ME_L5L6_L4D3PHI3X2_CM_L5L6_L4D3PHI3X2_wr_en;
wire [5:0] CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI3X2(
.data_in(ME_L5L6_L4D3PHI3X2_CM_L5L6_L4D3PHI3X2),
.enable(ME_L5L6_L4D3PHI3X2_CM_L5L6_L4D3PHI3X2_wr_en),
.number_out(CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3),
.start(ME_L5L6_L4D3PHI3X2_start),
.done(CM_L5L6_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D3PHI4X1_CM_L5L6_L4D3PHI4X1;
wire ME_L5L6_L4D3PHI4X1_CM_L5L6_L4D3PHI4X1_wr_en;
wire [5:0] CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI4X1(
.data_in(ME_L5L6_L4D3PHI4X1_CM_L5L6_L4D3PHI4X1),
.enable(ME_L5L6_L4D3PHI4X1_CM_L5L6_L4D3PHI4X1_wr_en),
.number_out(CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3),
.start(ME_L5L6_L4D3PHI4X1_start),
.done(CM_L5L6_L4D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D3PHI4X2_CM_L5L6_L4D3PHI4X2;
wire ME_L5L6_L4D3PHI4X2_CM_L5L6_L4D3PHI4X2_wr_en;
wire [5:0] CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3_number;
wire [8:0] CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3_read_add;
wire [11:0] CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3;
CandidateMatch  CM_L5L6_L4D3PHI4X2(
.data_in(ME_L5L6_L4D3PHI4X2_CM_L5L6_L4D3PHI4X2),
.enable(ME_L5L6_L4D3PHI4X2_CM_L5L6_L4D3PHI4X2_wr_en),
.number_out(CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3_number),
.read_add(CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3_read_add),
.data_out(CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3),
.start(ME_L5L6_L4D3PHI4X2_start),
.done(CM_L5L6_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L4D3_L5L6_AP_L5L6_L4D3;
wire PR_L4D3_L5L6_AP_L5L6_L4D3_wr_en;
wire [8:0] AP_L5L6_L4D3_MC_L5L6_L4D3_read_add;
wire [55:0] AP_L5L6_L4D3_MC_L5L6_L4D3;
AllProj #(1'b0,1'b0) AP_L5L6_L4D3(
.data_in(PR_L4D3_L5L6_AP_L5L6_L4D3),
.enable(PR_L4D3_L5L6_AP_L5L6_L4D3_wr_en),
.read_add(AP_L5L6_L4D3_MC_L5L6_L4D3_read_add),
.data_out(AP_L5L6_L4D3_MC_L5L6_L4D3),
.start(PR_L4D3_L5L6_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L4D3_AS_L4D3n2;
wire VMR_L4D3_AS_L4D3n2_wr_en;
wire [10:0] AS_L4D3n2_MC_L5L6_L4D3_read_add;
wire [35:0] AS_L4D3n2_MC_L5L6_L4D3;
AllStubs  AS_L4D3n2(
.data_in(VMR_L4D3_AS_L4D3n2),
.enable(VMR_L4D3_AS_L4D3n2_wr_en),
.read_add_MC(AS_L4D3n2_MC_L5L6_L4D3_read_add),
.data_out_MC(AS_L4D3n2_MC_L5L6_L4D3),
.start(VMR_L4D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D4PHI1X1_CM_L5L6_L4D4PHI1X1;
wire ME_L5L6_L4D4PHI1X1_CM_L5L6_L4D4PHI1X1_wr_en;
wire [5:0] CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI1X1(
.data_in(ME_L5L6_L4D4PHI1X1_CM_L5L6_L4D4PHI1X1),
.enable(ME_L5L6_L4D4PHI1X1_CM_L5L6_L4D4PHI1X1_wr_en),
.number_out(CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4),
.start(ME_L5L6_L4D4PHI1X1_start),
.done(CM_L5L6_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D4PHI1X2_CM_L5L6_L4D4PHI1X2;
wire ME_L5L6_L4D4PHI1X2_CM_L5L6_L4D4PHI1X2_wr_en;
wire [5:0] CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI1X2(
.data_in(ME_L5L6_L4D4PHI1X2_CM_L5L6_L4D4PHI1X2),
.enable(ME_L5L6_L4D4PHI1X2_CM_L5L6_L4D4PHI1X2_wr_en),
.number_out(CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4),
.start(ME_L5L6_L4D4PHI1X2_start),
.done(CM_L5L6_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D4PHI2X1_CM_L5L6_L4D4PHI2X1;
wire ME_L5L6_L4D4PHI2X1_CM_L5L6_L4D4PHI2X1_wr_en;
wire [5:0] CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI2X1(
.data_in(ME_L5L6_L4D4PHI2X1_CM_L5L6_L4D4PHI2X1),
.enable(ME_L5L6_L4D4PHI2X1_CM_L5L6_L4D4PHI2X1_wr_en),
.number_out(CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4),
.start(ME_L5L6_L4D4PHI2X1_start),
.done(CM_L5L6_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D4PHI2X2_CM_L5L6_L4D4PHI2X2;
wire ME_L5L6_L4D4PHI2X2_CM_L5L6_L4D4PHI2X2_wr_en;
wire [5:0] CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI2X2(
.data_in(ME_L5L6_L4D4PHI2X2_CM_L5L6_L4D4PHI2X2),
.enable(ME_L5L6_L4D4PHI2X2_CM_L5L6_L4D4PHI2X2_wr_en),
.number_out(CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4),
.start(ME_L5L6_L4D4PHI2X2_start),
.done(CM_L5L6_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D4PHI3X1_CM_L5L6_L4D4PHI3X1;
wire ME_L5L6_L4D4PHI3X1_CM_L5L6_L4D4PHI3X1_wr_en;
wire [5:0] CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI3X1(
.data_in(ME_L5L6_L4D4PHI3X1_CM_L5L6_L4D4PHI3X1),
.enable(ME_L5L6_L4D4PHI3X1_CM_L5L6_L4D4PHI3X1_wr_en),
.number_out(CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4),
.start(ME_L5L6_L4D4PHI3X1_start),
.done(CM_L5L6_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D4PHI3X2_CM_L5L6_L4D4PHI3X2;
wire ME_L5L6_L4D4PHI3X2_CM_L5L6_L4D4PHI3X2_wr_en;
wire [5:0] CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI3X2(
.data_in(ME_L5L6_L4D4PHI3X2_CM_L5L6_L4D4PHI3X2),
.enable(ME_L5L6_L4D4PHI3X2_CM_L5L6_L4D4PHI3X2_wr_en),
.number_out(CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4),
.start(ME_L5L6_L4D4PHI3X2_start),
.done(CM_L5L6_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D4PHI4X1_CM_L5L6_L4D4PHI4X1;
wire ME_L5L6_L4D4PHI4X1_CM_L5L6_L4D4PHI4X1_wr_en;
wire [5:0] CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI4X1(
.data_in(ME_L5L6_L4D4PHI4X1_CM_L5L6_L4D4PHI4X1),
.enable(ME_L5L6_L4D4PHI4X1_CM_L5L6_L4D4PHI4X1_wr_en),
.number_out(CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4),
.start(ME_L5L6_L4D4PHI4X1_start),
.done(CM_L5L6_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L5L6_L4D4PHI4X2_CM_L5L6_L4D4PHI4X2;
wire ME_L5L6_L4D4PHI4X2_CM_L5L6_L4D4PHI4X2_wr_en;
wire [5:0] CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4_number;
wire [8:0] CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4_read_add;
wire [11:0] CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4;
CandidateMatch  CM_L5L6_L4D4PHI4X2(
.data_in(ME_L5L6_L4D4PHI4X2_CM_L5L6_L4D4PHI4X2),
.enable(ME_L5L6_L4D4PHI4X2_CM_L5L6_L4D4PHI4X2_wr_en),
.number_out(CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4_number),
.read_add(CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4_read_add),
.data_out(CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4),
.start(ME_L5L6_L4D4PHI4X2_start),
.done(CM_L5L6_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L4D4_L5L6_AP_L5L6_L4D4;
wire PR_L4D4_L5L6_AP_L5L6_L4D4_wr_en;
wire [8:0] AP_L5L6_L4D4_MC_L5L6_L4D4_read_add;
wire [55:0] AP_L5L6_L4D4_MC_L5L6_L4D4;
AllProj #(1'b0,1'b0) AP_L5L6_L4D4(
.data_in(PR_L4D4_L5L6_AP_L5L6_L4D4),
.enable(PR_L4D4_L5L6_AP_L5L6_L4D4_wr_en),
.read_add(AP_L5L6_L4D4_MC_L5L6_L4D4_read_add),
.data_out(AP_L5L6_L4D4_MC_L5L6_L4D4),
.start(PR_L4D4_L5L6_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L4D4_AS_L4D4n3;
wire VMR_L4D4_AS_L4D4n3_wr_en;
wire [10:0] AS_L4D4n3_MC_L5L6_L4D4_read_add;
wire [35:0] AS_L4D4n3_MC_L5L6_L4D4;
AllStubs  AS_L4D4n3(
.data_in(VMR_L4D4_AS_L4D4n3),
.enable(VMR_L4D4_AS_L4D4n3_wr_en),
.read_add_MC(AS_L4D4n3_MC_L5L6_L4D4_read_add),
.data_out_MC(AS_L4D4n3_MC_L5L6_L4D4),
.start(VMR_L4D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D3PHI1X1_CM_L1L2_L3D3PHI1X1;
wire ME_L1L2_L3D3PHI1X1_CM_L1L2_L3D3PHI1X1_wr_en;
wire [5:0] CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI1X1(
.data_in(ME_L1L2_L3D3PHI1X1_CM_L1L2_L3D3PHI1X1),
.enable(ME_L1L2_L3D3PHI1X1_CM_L1L2_L3D3PHI1X1_wr_en),
.number_out(CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3),
.start(ME_L1L2_L3D3PHI1X1_start),
.done(CM_L1L2_L3D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D3PHI1X2_CM_L1L2_L3D3PHI1X2;
wire ME_L1L2_L3D3PHI1X2_CM_L1L2_L3D3PHI1X2_wr_en;
wire [5:0] CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI1X2(
.data_in(ME_L1L2_L3D3PHI1X2_CM_L1L2_L3D3PHI1X2),
.enable(ME_L1L2_L3D3PHI1X2_CM_L1L2_L3D3PHI1X2_wr_en),
.number_out(CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3),
.start(ME_L1L2_L3D3PHI1X2_start),
.done(CM_L1L2_L3D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D3PHI2X1_CM_L1L2_L3D3PHI2X1;
wire ME_L1L2_L3D3PHI2X1_CM_L1L2_L3D3PHI2X1_wr_en;
wire [5:0] CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI2X1(
.data_in(ME_L1L2_L3D3PHI2X1_CM_L1L2_L3D3PHI2X1),
.enable(ME_L1L2_L3D3PHI2X1_CM_L1L2_L3D3PHI2X1_wr_en),
.number_out(CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3),
.start(ME_L1L2_L3D3PHI2X1_start),
.done(CM_L1L2_L3D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D3PHI2X2_CM_L1L2_L3D3PHI2X2;
wire ME_L1L2_L3D3PHI2X2_CM_L1L2_L3D3PHI2X2_wr_en;
wire [5:0] CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI2X2(
.data_in(ME_L1L2_L3D3PHI2X2_CM_L1L2_L3D3PHI2X2),
.enable(ME_L1L2_L3D3PHI2X2_CM_L1L2_L3D3PHI2X2_wr_en),
.number_out(CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3),
.start(ME_L1L2_L3D3PHI2X2_start),
.done(CM_L1L2_L3D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D3PHI3X1_CM_L1L2_L3D3PHI3X1;
wire ME_L1L2_L3D3PHI3X1_CM_L1L2_L3D3PHI3X1_wr_en;
wire [5:0] CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI3X1(
.data_in(ME_L1L2_L3D3PHI3X1_CM_L1L2_L3D3PHI3X1),
.enable(ME_L1L2_L3D3PHI3X1_CM_L1L2_L3D3PHI3X1_wr_en),
.number_out(CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3),
.start(ME_L1L2_L3D3PHI3X1_start),
.done(CM_L1L2_L3D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D3PHI3X2_CM_L1L2_L3D3PHI3X2;
wire ME_L1L2_L3D3PHI3X2_CM_L1L2_L3D3PHI3X2_wr_en;
wire [5:0] CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3_number;
wire [8:0] CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3_read_add;
wire [11:0] CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3;
CandidateMatch  CM_L1L2_L3D3PHI3X2(
.data_in(ME_L1L2_L3D3PHI3X2_CM_L1L2_L3D3PHI3X2),
.enable(ME_L1L2_L3D3PHI3X2_CM_L1L2_L3D3PHI3X2_wr_en),
.number_out(CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3_number),
.read_add(CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3_read_add),
.data_out(CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3),
.start(ME_L1L2_L3D3PHI3X2_start),
.done(CM_L1L2_L3D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L3D3_L1L2_AP_L1L2_L3D3;
wire PR_L3D3_L1L2_AP_L1L2_L3D3_wr_en;
wire [8:0] AP_L1L2_L3D3_MC_L1L2_L3D3_read_add;
wire [55:0] AP_L1L2_L3D3_MC_L1L2_L3D3;
AllProj  AP_L1L2_L3D3(
.data_in(PR_L3D3_L1L2_AP_L1L2_L3D3),
.enable(PR_L3D3_L1L2_AP_L1L2_L3D3_wr_en),
.read_add(AP_L1L2_L3D3_MC_L1L2_L3D3_read_add),
.data_out(AP_L1L2_L3D3_MC_L1L2_L3D3),
.start(PR_L3D3_L1L2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L3D3_AS_L3D3n4;
wire VMR_L3D3_AS_L3D3n4_wr_en;
wire [10:0] AS_L3D3n4_MC_L1L2_L3D3_read_add;
wire [35:0] AS_L3D3n4_MC_L1L2_L3D3;
AllStubs  AS_L3D3n4(
.data_in(VMR_L3D3_AS_L3D3n4),
.enable(VMR_L3D3_AS_L3D3n4_wr_en),
.read_add_MC(AS_L3D3n4_MC_L1L2_L3D3_read_add),
.data_out_MC(AS_L3D3n4_MC_L1L2_L3D3),
.start(VMR_L3D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D4PHI1X1_CM_L1L2_L3D4PHI1X1;
wire ME_L1L2_L3D4PHI1X1_CM_L1L2_L3D4PHI1X1_wr_en;
wire [5:0] CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI1X1(
.data_in(ME_L1L2_L3D4PHI1X1_CM_L1L2_L3D4PHI1X1),
.enable(ME_L1L2_L3D4PHI1X1_CM_L1L2_L3D4PHI1X1_wr_en),
.number_out(CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4),
.start(ME_L1L2_L3D4PHI1X1_start),
.done(CM_L1L2_L3D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D4PHI1X2_CM_L1L2_L3D4PHI1X2;
wire ME_L1L2_L3D4PHI1X2_CM_L1L2_L3D4PHI1X2_wr_en;
wire [5:0] CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI1X2(
.data_in(ME_L1L2_L3D4PHI1X2_CM_L1L2_L3D4PHI1X2),
.enable(ME_L1L2_L3D4PHI1X2_CM_L1L2_L3D4PHI1X2_wr_en),
.number_out(CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4),
.start(ME_L1L2_L3D4PHI1X2_start),
.done(CM_L1L2_L3D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D4PHI2X1_CM_L1L2_L3D4PHI2X1;
wire ME_L1L2_L3D4PHI2X1_CM_L1L2_L3D4PHI2X1_wr_en;
wire [5:0] CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI2X1(
.data_in(ME_L1L2_L3D4PHI2X1_CM_L1L2_L3D4PHI2X1),
.enable(ME_L1L2_L3D4PHI2X1_CM_L1L2_L3D4PHI2X1_wr_en),
.number_out(CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4),
.start(ME_L1L2_L3D4PHI2X1_start),
.done(CM_L1L2_L3D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D4PHI2X2_CM_L1L2_L3D4PHI2X2;
wire ME_L1L2_L3D4PHI2X2_CM_L1L2_L3D4PHI2X2_wr_en;
wire [5:0] CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI2X2(
.data_in(ME_L1L2_L3D4PHI2X2_CM_L1L2_L3D4PHI2X2),
.enable(ME_L1L2_L3D4PHI2X2_CM_L1L2_L3D4PHI2X2_wr_en),
.number_out(CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4),
.start(ME_L1L2_L3D4PHI2X2_start),
.done(CM_L1L2_L3D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D4PHI3X1_CM_L1L2_L3D4PHI3X1;
wire ME_L1L2_L3D4PHI3X1_CM_L1L2_L3D4PHI3X1_wr_en;
wire [5:0] CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI3X1(
.data_in(ME_L1L2_L3D4PHI3X1_CM_L1L2_L3D4PHI3X1),
.enable(ME_L1L2_L3D4PHI3X1_CM_L1L2_L3D4PHI3X1_wr_en),
.number_out(CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4),
.start(ME_L1L2_L3D4PHI3X1_start),
.done(CM_L1L2_L3D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L3D4PHI3X2_CM_L1L2_L3D4PHI3X2;
wire ME_L1L2_L3D4PHI3X2_CM_L1L2_L3D4PHI3X2_wr_en;
wire [5:0] CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4_number;
wire [8:0] CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4_read_add;
wire [11:0] CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4;
CandidateMatch  CM_L1L2_L3D4PHI3X2(
.data_in(ME_L1L2_L3D4PHI3X2_CM_L1L2_L3D4PHI3X2),
.enable(ME_L1L2_L3D4PHI3X2_CM_L1L2_L3D4PHI3X2_wr_en),
.number_out(CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4_number),
.read_add(CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4_read_add),
.data_out(CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4),
.start(ME_L1L2_L3D4PHI3X2_start),
.done(CM_L1L2_L3D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L3D4_L1L2_AP_L1L2_L3D4;
wire PR_L3D4_L1L2_AP_L1L2_L3D4_wr_en;
wire [8:0] AP_L1L2_L3D4_MC_L1L2_L3D4_read_add;
wire [55:0] AP_L1L2_L3D4_MC_L1L2_L3D4;
AllProj  AP_L1L2_L3D4(
.data_in(PR_L3D4_L1L2_AP_L1L2_L3D4),
.enable(PR_L3D4_L1L2_AP_L1L2_L3D4_wr_en),
.read_add(AP_L1L2_L3D4_MC_L1L2_L3D4_read_add),
.data_out(AP_L1L2_L3D4_MC_L1L2_L3D4),
.start(PR_L3D4_L1L2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L3D4_AS_L3D4n3;
wire VMR_L3D4_AS_L3D4n3_wr_en;
wire [10:0] AS_L3D4n3_MC_L1L2_L3D4_read_add;
wire [35:0] AS_L3D4n3_MC_L1L2_L3D4;
AllStubs  AS_L3D4n3(
.data_in(VMR_L3D4_AS_L3D4n3),
.enable(VMR_L3D4_AS_L3D4n3_wr_en),
.read_add_MC(AS_L3D4n3_MC_L1L2_L3D4_read_add),
.data_out_MC(AS_L3D4n3_MC_L1L2_L3D4),
.start(VMR_L3D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D3PHI1X1_CM_L1L2_L4D3PHI1X1;
wire ME_L1L2_L4D3PHI1X1_CM_L1L2_L4D3PHI1X1_wr_en;
wire [5:0] CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI1X1(
.data_in(ME_L1L2_L4D3PHI1X1_CM_L1L2_L4D3PHI1X1),
.enable(ME_L1L2_L4D3PHI1X1_CM_L1L2_L4D3PHI1X1_wr_en),
.number_out(CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3),
.start(ME_L1L2_L4D3PHI1X1_start),
.done(CM_L1L2_L4D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D3PHI1X2_CM_L1L2_L4D3PHI1X2;
wire ME_L1L2_L4D3PHI1X2_CM_L1L2_L4D3PHI1X2_wr_en;
wire [5:0] CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI1X2(
.data_in(ME_L1L2_L4D3PHI1X2_CM_L1L2_L4D3PHI1X2),
.enable(ME_L1L2_L4D3PHI1X2_CM_L1L2_L4D3PHI1X2_wr_en),
.number_out(CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3),
.start(ME_L1L2_L4D3PHI1X2_start),
.done(CM_L1L2_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D3PHI2X1_CM_L1L2_L4D3PHI2X1;
wire ME_L1L2_L4D3PHI2X1_CM_L1L2_L4D3PHI2X1_wr_en;
wire [5:0] CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI2X1(
.data_in(ME_L1L2_L4D3PHI2X1_CM_L1L2_L4D3PHI2X1),
.enable(ME_L1L2_L4D3PHI2X1_CM_L1L2_L4D3PHI2X1_wr_en),
.number_out(CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3),
.start(ME_L1L2_L4D3PHI2X1_start),
.done(CM_L1L2_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D3PHI2X2_CM_L1L2_L4D3PHI2X2;
wire ME_L1L2_L4D3PHI2X2_CM_L1L2_L4D3PHI2X2_wr_en;
wire [5:0] CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI2X2(
.data_in(ME_L1L2_L4D3PHI2X2_CM_L1L2_L4D3PHI2X2),
.enable(ME_L1L2_L4D3PHI2X2_CM_L1L2_L4D3PHI2X2_wr_en),
.number_out(CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3),
.start(ME_L1L2_L4D3PHI2X2_start),
.done(CM_L1L2_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D3PHI3X1_CM_L1L2_L4D3PHI3X1;
wire ME_L1L2_L4D3PHI3X1_CM_L1L2_L4D3PHI3X1_wr_en;
wire [5:0] CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI3X1(
.data_in(ME_L1L2_L4D3PHI3X1_CM_L1L2_L4D3PHI3X1),
.enable(ME_L1L2_L4D3PHI3X1_CM_L1L2_L4D3PHI3X1_wr_en),
.number_out(CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3),
.start(ME_L1L2_L4D3PHI3X1_start),
.done(CM_L1L2_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D3PHI3X2_CM_L1L2_L4D3PHI3X2;
wire ME_L1L2_L4D3PHI3X2_CM_L1L2_L4D3PHI3X2_wr_en;
wire [5:0] CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI3X2(
.data_in(ME_L1L2_L4D3PHI3X2_CM_L1L2_L4D3PHI3X2),
.enable(ME_L1L2_L4D3PHI3X2_CM_L1L2_L4D3PHI3X2_wr_en),
.number_out(CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3),
.start(ME_L1L2_L4D3PHI3X2_start),
.done(CM_L1L2_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D3PHI4X1_CM_L1L2_L4D3PHI4X1;
wire ME_L1L2_L4D3PHI4X1_CM_L1L2_L4D3PHI4X1_wr_en;
wire [5:0] CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI4X1(
.data_in(ME_L1L2_L4D3PHI4X1_CM_L1L2_L4D3PHI4X1),
.enable(ME_L1L2_L4D3PHI4X1_CM_L1L2_L4D3PHI4X1_wr_en),
.number_out(CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3),
.start(ME_L1L2_L4D3PHI4X1_start),
.done(CM_L1L2_L4D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D3PHI4X2_CM_L1L2_L4D3PHI4X2;
wire ME_L1L2_L4D3PHI4X2_CM_L1L2_L4D3PHI4X2_wr_en;
wire [5:0] CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3_number;
wire [8:0] CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3_read_add;
wire [11:0] CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3;
CandidateMatch  CM_L1L2_L4D3PHI4X2(
.data_in(ME_L1L2_L4D3PHI4X2_CM_L1L2_L4D3PHI4X2),
.enable(ME_L1L2_L4D3PHI4X2_CM_L1L2_L4D3PHI4X2_wr_en),
.number_out(CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3_number),
.read_add(CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3_read_add),
.data_out(CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3),
.start(ME_L1L2_L4D3PHI4X2_start),
.done(CM_L1L2_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L4D3_L1L2_AP_L1L2_L4D3;
wire PR_L4D3_L1L2_AP_L1L2_L4D3_wr_en;
wire [8:0] AP_L1L2_L4D3_MC_L1L2_L4D3_read_add;
wire [55:0] AP_L1L2_L4D3_MC_L1L2_L4D3;
AllProj #(1'b0,1'b0) AP_L1L2_L4D3(
.data_in(PR_L4D3_L1L2_AP_L1L2_L4D3),
.enable(PR_L4D3_L1L2_AP_L1L2_L4D3_wr_en),
.read_add(AP_L1L2_L4D3_MC_L1L2_L4D3_read_add),
.data_out(AP_L1L2_L4D3_MC_L1L2_L4D3),
.start(PR_L4D3_L1L2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L4D3_AS_L4D3n3;
wire VMR_L4D3_AS_L4D3n3_wr_en;
wire [10:0] AS_L4D3n3_MC_L1L2_L4D3_read_add;
wire [35:0] AS_L4D3n3_MC_L1L2_L4D3;
AllStubs  AS_L4D3n3(
.data_in(VMR_L4D3_AS_L4D3n3),
.enable(VMR_L4D3_AS_L4D3n3_wr_en),
.read_add_MC(AS_L4D3n3_MC_L1L2_L4D3_read_add),
.data_out_MC(AS_L4D3n3_MC_L1L2_L4D3),
.start(VMR_L4D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D4PHI1X1_CM_L1L2_L4D4PHI1X1;
wire ME_L1L2_L4D4PHI1X1_CM_L1L2_L4D4PHI1X1_wr_en;
wire [5:0] CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI1X1(
.data_in(ME_L1L2_L4D4PHI1X1_CM_L1L2_L4D4PHI1X1),
.enable(ME_L1L2_L4D4PHI1X1_CM_L1L2_L4D4PHI1X1_wr_en),
.number_out(CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4),
.start(ME_L1L2_L4D4PHI1X1_start),
.done(CM_L1L2_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D4PHI1X2_CM_L1L2_L4D4PHI1X2;
wire ME_L1L2_L4D4PHI1X2_CM_L1L2_L4D4PHI1X2_wr_en;
wire [5:0] CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI1X2(
.data_in(ME_L1L2_L4D4PHI1X2_CM_L1L2_L4D4PHI1X2),
.enable(ME_L1L2_L4D4PHI1X2_CM_L1L2_L4D4PHI1X2_wr_en),
.number_out(CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4),
.start(ME_L1L2_L4D4PHI1X2_start),
.done(CM_L1L2_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D4PHI2X1_CM_L1L2_L4D4PHI2X1;
wire ME_L1L2_L4D4PHI2X1_CM_L1L2_L4D4PHI2X1_wr_en;
wire [5:0] CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI2X1(
.data_in(ME_L1L2_L4D4PHI2X1_CM_L1L2_L4D4PHI2X1),
.enable(ME_L1L2_L4D4PHI2X1_CM_L1L2_L4D4PHI2X1_wr_en),
.number_out(CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4),
.start(ME_L1L2_L4D4PHI2X1_start),
.done(CM_L1L2_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D4PHI2X2_CM_L1L2_L4D4PHI2X2;
wire ME_L1L2_L4D4PHI2X2_CM_L1L2_L4D4PHI2X2_wr_en;
wire [5:0] CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI2X2(
.data_in(ME_L1L2_L4D4PHI2X2_CM_L1L2_L4D4PHI2X2),
.enable(ME_L1L2_L4D4PHI2X2_CM_L1L2_L4D4PHI2X2_wr_en),
.number_out(CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4),
.start(ME_L1L2_L4D4PHI2X2_start),
.done(CM_L1L2_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D4PHI3X1_CM_L1L2_L4D4PHI3X1;
wire ME_L1L2_L4D4PHI3X1_CM_L1L2_L4D4PHI3X1_wr_en;
wire [5:0] CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI3X1(
.data_in(ME_L1L2_L4D4PHI3X1_CM_L1L2_L4D4PHI3X1),
.enable(ME_L1L2_L4D4PHI3X1_CM_L1L2_L4D4PHI3X1_wr_en),
.number_out(CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4),
.start(ME_L1L2_L4D4PHI3X1_start),
.done(CM_L1L2_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D4PHI3X2_CM_L1L2_L4D4PHI3X2;
wire ME_L1L2_L4D4PHI3X2_CM_L1L2_L4D4PHI3X2_wr_en;
wire [5:0] CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI3X2(
.data_in(ME_L1L2_L4D4PHI3X2_CM_L1L2_L4D4PHI3X2),
.enable(ME_L1L2_L4D4PHI3X2_CM_L1L2_L4D4PHI3X2_wr_en),
.number_out(CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4),
.start(ME_L1L2_L4D4PHI3X2_start),
.done(CM_L1L2_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D4PHI4X1_CM_L1L2_L4D4PHI4X1;
wire ME_L1L2_L4D4PHI4X1_CM_L1L2_L4D4PHI4X1_wr_en;
wire [5:0] CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI4X1(
.data_in(ME_L1L2_L4D4PHI4X1_CM_L1L2_L4D4PHI4X1),
.enable(ME_L1L2_L4D4PHI4X1_CM_L1L2_L4D4PHI4X1_wr_en),
.number_out(CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4),
.start(ME_L1L2_L4D4PHI4X1_start),
.done(CM_L1L2_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L4D4PHI4X2_CM_L1L2_L4D4PHI4X2;
wire ME_L1L2_L4D4PHI4X2_CM_L1L2_L4D4PHI4X2_wr_en;
wire [5:0] CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4_number;
wire [8:0] CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4_read_add;
wire [11:0] CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4;
CandidateMatch  CM_L1L2_L4D4PHI4X2(
.data_in(ME_L1L2_L4D4PHI4X2_CM_L1L2_L4D4PHI4X2),
.enable(ME_L1L2_L4D4PHI4X2_CM_L1L2_L4D4PHI4X2_wr_en),
.number_out(CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4_number),
.read_add(CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4_read_add),
.data_out(CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4),
.start(ME_L1L2_L4D4PHI4X2_start),
.done(CM_L1L2_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L4D4_L1L2_AP_L1L2_L4D4;
wire PR_L4D4_L1L2_AP_L1L2_L4D4_wr_en;
wire [8:0] AP_L1L2_L4D4_MC_L1L2_L4D4_read_add;
wire [55:0] AP_L1L2_L4D4_MC_L1L2_L4D4;
AllProj #(1'b0,1'b0) AP_L1L2_L4D4(
.data_in(PR_L4D4_L1L2_AP_L1L2_L4D4),
.enable(PR_L4D4_L1L2_AP_L1L2_L4D4_wr_en),
.read_add(AP_L1L2_L4D4_MC_L1L2_L4D4_read_add),
.data_out(AP_L1L2_L4D4_MC_L1L2_L4D4),
.start(PR_L4D4_L1L2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L4D4_AS_L4D4n4;
wire VMR_L4D4_AS_L4D4n4_wr_en;
wire [10:0] AS_L4D4n4_MC_L1L2_L4D4_read_add;
wire [35:0] AS_L4D4n4_MC_L1L2_L4D4;
AllStubs  AS_L4D4n4(
.data_in(VMR_L4D4_AS_L4D4n4),
.enable(VMR_L4D4_AS_L4D4n4_wr_en),
.read_add_MC(AS_L4D4n4_MC_L1L2_L4D4_read_add),
.data_out_MC(AS_L4D4n4_MC_L1L2_L4D4),
.start(VMR_L4D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D3PHI1X1_CM_L1L2_L5D3PHI1X1;
wire ME_L1L2_L5D3PHI1X1_CM_L1L2_L5D3PHI1X1_wr_en;
wire [5:0] CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI1X1(
.data_in(ME_L1L2_L5D3PHI1X1_CM_L1L2_L5D3PHI1X1),
.enable(ME_L1L2_L5D3PHI1X1_CM_L1L2_L5D3PHI1X1_wr_en),
.number_out(CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3),
.start(ME_L1L2_L5D3PHI1X1_start),
.done(CM_L1L2_L5D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D3PHI1X2_CM_L1L2_L5D3PHI1X2;
wire ME_L1L2_L5D3PHI1X2_CM_L1L2_L5D3PHI1X2_wr_en;
wire [5:0] CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI1X2(
.data_in(ME_L1L2_L5D3PHI1X2_CM_L1L2_L5D3PHI1X2),
.enable(ME_L1L2_L5D3PHI1X2_CM_L1L2_L5D3PHI1X2_wr_en),
.number_out(CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3),
.start(ME_L1L2_L5D3PHI1X2_start),
.done(CM_L1L2_L5D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D3PHI2X1_CM_L1L2_L5D3PHI2X1;
wire ME_L1L2_L5D3PHI2X1_CM_L1L2_L5D3PHI2X1_wr_en;
wire [5:0] CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI2X1(
.data_in(ME_L1L2_L5D3PHI2X1_CM_L1L2_L5D3PHI2X1),
.enable(ME_L1L2_L5D3PHI2X1_CM_L1L2_L5D3PHI2X1_wr_en),
.number_out(CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3),
.start(ME_L1L2_L5D3PHI2X1_start),
.done(CM_L1L2_L5D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D3PHI2X2_CM_L1L2_L5D3PHI2X2;
wire ME_L1L2_L5D3PHI2X2_CM_L1L2_L5D3PHI2X2_wr_en;
wire [5:0] CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI2X2(
.data_in(ME_L1L2_L5D3PHI2X2_CM_L1L2_L5D3PHI2X2),
.enable(ME_L1L2_L5D3PHI2X2_CM_L1L2_L5D3PHI2X2_wr_en),
.number_out(CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3),
.start(ME_L1L2_L5D3PHI2X2_start),
.done(CM_L1L2_L5D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D3PHI3X1_CM_L1L2_L5D3PHI3X1;
wire ME_L1L2_L5D3PHI3X1_CM_L1L2_L5D3PHI3X1_wr_en;
wire [5:0] CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI3X1(
.data_in(ME_L1L2_L5D3PHI3X1_CM_L1L2_L5D3PHI3X1),
.enable(ME_L1L2_L5D3PHI3X1_CM_L1L2_L5D3PHI3X1_wr_en),
.number_out(CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3),
.start(ME_L1L2_L5D3PHI3X1_start),
.done(CM_L1L2_L5D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D3PHI3X2_CM_L1L2_L5D3PHI3X2;
wire ME_L1L2_L5D3PHI3X2_CM_L1L2_L5D3PHI3X2_wr_en;
wire [5:0] CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3_number;
wire [8:0] CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3_read_add;
wire [11:0] CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3;
CandidateMatch  CM_L1L2_L5D3PHI3X2(
.data_in(ME_L1L2_L5D3PHI3X2_CM_L1L2_L5D3PHI3X2),
.enable(ME_L1L2_L5D3PHI3X2_CM_L1L2_L5D3PHI3X2_wr_en),
.number_out(CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3_number),
.read_add(CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3_read_add),
.data_out(CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3),
.start(ME_L1L2_L5D3PHI3X2_start),
.done(CM_L1L2_L5D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L5D3_L1L2_AP_L1L2_L5D3;
wire PR_L5D3_L1L2_AP_L1L2_L5D3_wr_en;
wire [8:0] AP_L1L2_L5D3_MC_L1L2_L5D3_read_add;
wire [55:0] AP_L1L2_L5D3_MC_L1L2_L5D3;
AllProj #(1'b0,1'b0) AP_L1L2_L5D3(
.data_in(PR_L5D3_L1L2_AP_L1L2_L5D3),
.enable(PR_L5D3_L1L2_AP_L1L2_L5D3_wr_en),
.read_add(AP_L1L2_L5D3_MC_L1L2_L5D3_read_add),
.data_out(AP_L1L2_L5D3_MC_L1L2_L5D3),
.start(PR_L5D3_L1L2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L5D3_AS_L5D3n4;
wire VMR_L5D3_AS_L5D3n4_wr_en;
wire [10:0] AS_L5D3n4_MC_L1L2_L5D3_read_add;
wire [35:0] AS_L5D3n4_MC_L1L2_L5D3;
AllStubs  AS_L5D3n4(
.data_in(VMR_L5D3_AS_L5D3n4),
.enable(VMR_L5D3_AS_L5D3n4_wr_en),
.read_add_MC(AS_L5D3n4_MC_L1L2_L5D3_read_add),
.data_out_MC(AS_L5D3n4_MC_L1L2_L5D3),
.start(VMR_L5D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D4PHI1X1_CM_L1L2_L5D4PHI1X1;
wire ME_L1L2_L5D4PHI1X1_CM_L1L2_L5D4PHI1X1_wr_en;
wire [5:0] CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI1X1(
.data_in(ME_L1L2_L5D4PHI1X1_CM_L1L2_L5D4PHI1X1),
.enable(ME_L1L2_L5D4PHI1X1_CM_L1L2_L5D4PHI1X1_wr_en),
.number_out(CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4),
.start(ME_L1L2_L5D4PHI1X1_start),
.done(CM_L1L2_L5D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D4PHI1X2_CM_L1L2_L5D4PHI1X2;
wire ME_L1L2_L5D4PHI1X2_CM_L1L2_L5D4PHI1X2_wr_en;
wire [5:0] CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI1X2(
.data_in(ME_L1L2_L5D4PHI1X2_CM_L1L2_L5D4PHI1X2),
.enable(ME_L1L2_L5D4PHI1X2_CM_L1L2_L5D4PHI1X2_wr_en),
.number_out(CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4),
.start(ME_L1L2_L5D4PHI1X2_start),
.done(CM_L1L2_L5D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D4PHI2X1_CM_L1L2_L5D4PHI2X1;
wire ME_L1L2_L5D4PHI2X1_CM_L1L2_L5D4PHI2X1_wr_en;
wire [5:0] CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI2X1(
.data_in(ME_L1L2_L5D4PHI2X1_CM_L1L2_L5D4PHI2X1),
.enable(ME_L1L2_L5D4PHI2X1_CM_L1L2_L5D4PHI2X1_wr_en),
.number_out(CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4),
.start(ME_L1L2_L5D4PHI2X1_start),
.done(CM_L1L2_L5D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D4PHI2X2_CM_L1L2_L5D4PHI2X2;
wire ME_L1L2_L5D4PHI2X2_CM_L1L2_L5D4PHI2X2_wr_en;
wire [5:0] CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI2X2(
.data_in(ME_L1L2_L5D4PHI2X2_CM_L1L2_L5D4PHI2X2),
.enable(ME_L1L2_L5D4PHI2X2_CM_L1L2_L5D4PHI2X2_wr_en),
.number_out(CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4),
.start(ME_L1L2_L5D4PHI2X2_start),
.done(CM_L1L2_L5D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D4PHI3X1_CM_L1L2_L5D4PHI3X1;
wire ME_L1L2_L5D4PHI3X1_CM_L1L2_L5D4PHI3X1_wr_en;
wire [5:0] CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI3X1(
.data_in(ME_L1L2_L5D4PHI3X1_CM_L1L2_L5D4PHI3X1),
.enable(ME_L1L2_L5D4PHI3X1_CM_L1L2_L5D4PHI3X1_wr_en),
.number_out(CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4),
.start(ME_L1L2_L5D4PHI3X1_start),
.done(CM_L1L2_L5D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L5D4PHI3X2_CM_L1L2_L5D4PHI3X2;
wire ME_L1L2_L5D4PHI3X2_CM_L1L2_L5D4PHI3X2_wr_en;
wire [5:0] CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4_number;
wire [8:0] CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4_read_add;
wire [11:0] CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4;
CandidateMatch  CM_L1L2_L5D4PHI3X2(
.data_in(ME_L1L2_L5D4PHI3X2_CM_L1L2_L5D4PHI3X2),
.enable(ME_L1L2_L5D4PHI3X2_CM_L1L2_L5D4PHI3X2_wr_en),
.number_out(CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4_number),
.read_add(CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4_read_add),
.data_out(CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4),
.start(ME_L1L2_L5D4PHI3X2_start),
.done(CM_L1L2_L5D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L5D4_L1L2_AP_L1L2_L5D4;
wire PR_L5D4_L1L2_AP_L1L2_L5D4_wr_en;
wire [8:0] AP_L1L2_L5D4_MC_L1L2_L5D4_read_add;
wire [55:0] AP_L1L2_L5D4_MC_L1L2_L5D4;
AllProj #(1'b0,1'b0) AP_L1L2_L5D4(
.data_in(PR_L5D4_L1L2_AP_L1L2_L5D4),
.enable(PR_L5D4_L1L2_AP_L1L2_L5D4_wr_en),
.read_add(AP_L1L2_L5D4_MC_L1L2_L5D4_read_add),
.data_out(AP_L1L2_L5D4_MC_L1L2_L5D4),
.start(PR_L5D4_L1L2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L5D4_AS_L5D4n3;
wire VMR_L5D4_AS_L5D4n3_wr_en;
wire [10:0] AS_L5D4n3_MC_L1L2_L5D4_read_add;
wire [35:0] AS_L5D4n3_MC_L1L2_L5D4;
AllStubs  AS_L5D4n3(
.data_in(VMR_L5D4_AS_L5D4n3),
.enable(VMR_L5D4_AS_L5D4n3_wr_en),
.read_add_MC(AS_L5D4n3_MC_L1L2_L5D4_read_add),
.data_out_MC(AS_L5D4n3_MC_L1L2_L5D4),
.start(VMR_L5D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D3PHI1X1_CM_L1L2_L6D3PHI1X1;
wire ME_L1L2_L6D3PHI1X1_CM_L1L2_L6D3PHI1X1_wr_en;
wire [5:0] CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI1X1(
.data_in(ME_L1L2_L6D3PHI1X1_CM_L1L2_L6D3PHI1X1),
.enable(ME_L1L2_L6D3PHI1X1_CM_L1L2_L6D3PHI1X1_wr_en),
.number_out(CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3),
.start(ME_L1L2_L6D3PHI1X1_start),
.done(CM_L1L2_L6D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D3PHI1X2_CM_L1L2_L6D3PHI1X2;
wire ME_L1L2_L6D3PHI1X2_CM_L1L2_L6D3PHI1X2_wr_en;
wire [5:0] CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI1X2(
.data_in(ME_L1L2_L6D3PHI1X2_CM_L1L2_L6D3PHI1X2),
.enable(ME_L1L2_L6D3PHI1X2_CM_L1L2_L6D3PHI1X2_wr_en),
.number_out(CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3),
.start(ME_L1L2_L6D3PHI1X2_start),
.done(CM_L1L2_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D3PHI2X1_CM_L1L2_L6D3PHI2X1;
wire ME_L1L2_L6D3PHI2X1_CM_L1L2_L6D3PHI2X1_wr_en;
wire [5:0] CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI2X1(
.data_in(ME_L1L2_L6D3PHI2X1_CM_L1L2_L6D3PHI2X1),
.enable(ME_L1L2_L6D3PHI2X1_CM_L1L2_L6D3PHI2X1_wr_en),
.number_out(CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3),
.start(ME_L1L2_L6D3PHI2X1_start),
.done(CM_L1L2_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D3PHI2X2_CM_L1L2_L6D3PHI2X2;
wire ME_L1L2_L6D3PHI2X2_CM_L1L2_L6D3PHI2X2_wr_en;
wire [5:0] CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI2X2(
.data_in(ME_L1L2_L6D3PHI2X2_CM_L1L2_L6D3PHI2X2),
.enable(ME_L1L2_L6D3PHI2X2_CM_L1L2_L6D3PHI2X2_wr_en),
.number_out(CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3),
.start(ME_L1L2_L6D3PHI2X2_start),
.done(CM_L1L2_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D3PHI3X1_CM_L1L2_L6D3PHI3X1;
wire ME_L1L2_L6D3PHI3X1_CM_L1L2_L6D3PHI3X1_wr_en;
wire [5:0] CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI3X1(
.data_in(ME_L1L2_L6D3PHI3X1_CM_L1L2_L6D3PHI3X1),
.enable(ME_L1L2_L6D3PHI3X1_CM_L1L2_L6D3PHI3X1_wr_en),
.number_out(CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3),
.start(ME_L1L2_L6D3PHI3X1_start),
.done(CM_L1L2_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D3PHI3X2_CM_L1L2_L6D3PHI3X2;
wire ME_L1L2_L6D3PHI3X2_CM_L1L2_L6D3PHI3X2_wr_en;
wire [5:0] CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI3X2(
.data_in(ME_L1L2_L6D3PHI3X2_CM_L1L2_L6D3PHI3X2),
.enable(ME_L1L2_L6D3PHI3X2_CM_L1L2_L6D3PHI3X2_wr_en),
.number_out(CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3),
.start(ME_L1L2_L6D3PHI3X2_start),
.done(CM_L1L2_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D3PHI4X1_CM_L1L2_L6D3PHI4X1;
wire ME_L1L2_L6D3PHI4X1_CM_L1L2_L6D3PHI4X1_wr_en;
wire [5:0] CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI4X1(
.data_in(ME_L1L2_L6D3PHI4X1_CM_L1L2_L6D3PHI4X1),
.enable(ME_L1L2_L6D3PHI4X1_CM_L1L2_L6D3PHI4X1_wr_en),
.number_out(CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3),
.start(ME_L1L2_L6D3PHI4X1_start),
.done(CM_L1L2_L6D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D3PHI4X2_CM_L1L2_L6D3PHI4X2;
wire ME_L1L2_L6D3PHI4X2_CM_L1L2_L6D3PHI4X2_wr_en;
wire [5:0] CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3_number;
wire [8:0] CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3_read_add;
wire [11:0] CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3;
CandidateMatch  CM_L1L2_L6D3PHI4X2(
.data_in(ME_L1L2_L6D3PHI4X2_CM_L1L2_L6D3PHI4X2),
.enable(ME_L1L2_L6D3PHI4X2_CM_L1L2_L6D3PHI4X2_wr_en),
.number_out(CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3_number),
.read_add(CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3_read_add),
.data_out(CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3),
.start(ME_L1L2_L6D3PHI4X2_start),
.done(CM_L1L2_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L6D3_L1L2_AP_L1L2_L6D3;
wire PR_L6D3_L1L2_AP_L1L2_L6D3_wr_en;
wire [8:0] AP_L1L2_L6D3_MC_L1L2_L6D3_read_add;
wire [55:0] AP_L1L2_L6D3_MC_L1L2_L6D3;
AllProj #(1'b0,1'b0) AP_L1L2_L6D3(
.data_in(PR_L6D3_L1L2_AP_L1L2_L6D3),
.enable(PR_L6D3_L1L2_AP_L1L2_L6D3_wr_en),
.read_add(AP_L1L2_L6D3_MC_L1L2_L6D3_read_add),
.data_out(AP_L1L2_L6D3_MC_L1L2_L6D3),
.start(PR_L6D3_L1L2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L6D3_AS_L6D3n3;
wire VMR_L6D3_AS_L6D3n3_wr_en;
wire [10:0] AS_L6D3n3_MC_L1L2_L6D3_read_add;
wire [35:0] AS_L6D3n3_MC_L1L2_L6D3;
AllStubs  AS_L6D3n3(
.data_in(VMR_L6D3_AS_L6D3n3),
.enable(VMR_L6D3_AS_L6D3n3_wr_en),
.read_add_MC(AS_L6D3n3_MC_L1L2_L6D3_read_add),
.data_out_MC(AS_L6D3n3_MC_L1L2_L6D3),
.start(VMR_L6D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D4PHI1X1_CM_L1L2_L6D4PHI1X1;
wire ME_L1L2_L6D4PHI1X1_CM_L1L2_L6D4PHI1X1_wr_en;
wire [5:0] CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI1X1(
.data_in(ME_L1L2_L6D4PHI1X1_CM_L1L2_L6D4PHI1X1),
.enable(ME_L1L2_L6D4PHI1X1_CM_L1L2_L6D4PHI1X1_wr_en),
.number_out(CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4),
.start(ME_L1L2_L6D4PHI1X1_start),
.done(CM_L1L2_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D4PHI1X2_CM_L1L2_L6D4PHI1X2;
wire ME_L1L2_L6D4PHI1X2_CM_L1L2_L6D4PHI1X2_wr_en;
wire [5:0] CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI1X2(
.data_in(ME_L1L2_L6D4PHI1X2_CM_L1L2_L6D4PHI1X2),
.enable(ME_L1L2_L6D4PHI1X2_CM_L1L2_L6D4PHI1X2_wr_en),
.number_out(CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4),
.start(ME_L1L2_L6D4PHI1X2_start),
.done(CM_L1L2_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D4PHI2X1_CM_L1L2_L6D4PHI2X1;
wire ME_L1L2_L6D4PHI2X1_CM_L1L2_L6D4PHI2X1_wr_en;
wire [5:0] CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI2X1(
.data_in(ME_L1L2_L6D4PHI2X1_CM_L1L2_L6D4PHI2X1),
.enable(ME_L1L2_L6D4PHI2X1_CM_L1L2_L6D4PHI2X1_wr_en),
.number_out(CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4),
.start(ME_L1L2_L6D4PHI2X1_start),
.done(CM_L1L2_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D4PHI2X2_CM_L1L2_L6D4PHI2X2;
wire ME_L1L2_L6D4PHI2X2_CM_L1L2_L6D4PHI2X2_wr_en;
wire [5:0] CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI2X2(
.data_in(ME_L1L2_L6D4PHI2X2_CM_L1L2_L6D4PHI2X2),
.enable(ME_L1L2_L6D4PHI2X2_CM_L1L2_L6D4PHI2X2_wr_en),
.number_out(CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4),
.start(ME_L1L2_L6D4PHI2X2_start),
.done(CM_L1L2_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D4PHI3X1_CM_L1L2_L6D4PHI3X1;
wire ME_L1L2_L6D4PHI3X1_CM_L1L2_L6D4PHI3X1_wr_en;
wire [5:0] CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI3X1(
.data_in(ME_L1L2_L6D4PHI3X1_CM_L1L2_L6D4PHI3X1),
.enable(ME_L1L2_L6D4PHI3X1_CM_L1L2_L6D4PHI3X1_wr_en),
.number_out(CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4),
.start(ME_L1L2_L6D4PHI3X1_start),
.done(CM_L1L2_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D4PHI3X2_CM_L1L2_L6D4PHI3X2;
wire ME_L1L2_L6D4PHI3X2_CM_L1L2_L6D4PHI3X2_wr_en;
wire [5:0] CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI3X2(
.data_in(ME_L1L2_L6D4PHI3X2_CM_L1L2_L6D4PHI3X2),
.enable(ME_L1L2_L6D4PHI3X2_CM_L1L2_L6D4PHI3X2_wr_en),
.number_out(CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4),
.start(ME_L1L2_L6D4PHI3X2_start),
.done(CM_L1L2_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D4PHI4X1_CM_L1L2_L6D4PHI4X1;
wire ME_L1L2_L6D4PHI4X1_CM_L1L2_L6D4PHI4X1_wr_en;
wire [5:0] CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI4X1(
.data_in(ME_L1L2_L6D4PHI4X1_CM_L1L2_L6D4PHI4X1),
.enable(ME_L1L2_L6D4PHI4X1_CM_L1L2_L6D4PHI4X1_wr_en),
.number_out(CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4),
.start(ME_L1L2_L6D4PHI4X1_start),
.done(CM_L1L2_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [11:0] ME_L1L2_L6D4PHI4X2_CM_L1L2_L6D4PHI4X2;
wire ME_L1L2_L6D4PHI4X2_CM_L1L2_L6D4PHI4X2_wr_en;
wire [5:0] CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4_number;
wire [8:0] CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4_read_add;
wire [11:0] CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4;
CandidateMatch  CM_L1L2_L6D4PHI4X2(
.data_in(ME_L1L2_L6D4PHI4X2_CM_L1L2_L6D4PHI4X2),
.enable(ME_L1L2_L6D4PHI4X2_CM_L1L2_L6D4PHI4X2_wr_en),
.number_out(CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4_number),
.read_add(CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4_read_add),
.data_out(CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4),
.start(ME_L1L2_L6D4PHI4X2_start),
.done(CM_L1L2_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [55:0] PR_L6D4_L1L2_AP_L1L2_L6D4;
wire PR_L6D4_L1L2_AP_L1L2_L6D4_wr_en;
wire [8:0] AP_L1L2_L6D4_MC_L1L2_L6D4_read_add;
wire [55:0] AP_L1L2_L6D4_MC_L1L2_L6D4;
AllProj #(1'b0,1'b0) AP_L1L2_L6D4(
.data_in(PR_L6D4_L1L2_AP_L1L2_L6D4),
.enable(PR_L6D4_L1L2_AP_L1L2_L6D4_wr_en),
.read_add(AP_L1L2_L6D4_MC_L1L2_L6D4_read_add),
.data_out(AP_L1L2_L6D4_MC_L1L2_L6D4),
.start(PR_L6D4_L1L2_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [35:0] VMR_L6D4_AS_L6D4n4;
wire VMR_L6D4_AS_L6D4n4_wr_en;
wire [10:0] AS_L6D4n4_MC_L1L2_L6D4_read_add;
wire [35:0] AS_L6D4n4_MC_L1L2_L6D4;
AllStubs  AS_L6D4n4(
.data_in(VMR_L6D4_AS_L6D4n4),
.enable(VMR_L6D4_AS_L6D4n4_wr_en),
.read_add_MC(AS_L6D4n4_MC_L1L2_L6D4_read_add),
.data_out_MC(AS_L6D4n4_MC_L1L2_L6D4),
.start(VMR_L6D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus;
wire MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus_wr_en;
wire [5:0] FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L1L2_L3D3_ToMinus_MT_Layr_Minus;
wire FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L1L2_L3D3_ToMinus(
.data_in(MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus),
.enable(MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus_wr_en),
.number_out(FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L1L2_L3D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L1L2_L3D3_start),
.done(FM_L1L2_L3D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus;
wire MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus_wr_en;
wire [5:0] FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L1L2_L4D3_ToMinus_MT_Layr_Minus;
wire FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L1L2_L4D3_ToMinus(
.data_in(MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus),
.enable(MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus_wr_en),
.number_out(FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L1L2_L4D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L1L2_L4D3_start),
.done(FM_L1L2_L4D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus;
wire MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus_wr_en;
wire [5:0] FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L1L2_L5D3_ToMinus_MT_Layr_Minus;
wire FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L1L2_L5D3_ToMinus(
.data_in(MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus),
.enable(MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus_wr_en),
.number_out(FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L1L2_L5D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L1L2_L5D3_start),
.done(FM_L1L2_L5D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus;
wire MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus_wr_en;
wire [5:0] FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L1L2_L6D3_ToMinus_MT_Layr_Minus;
wire FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L1L2_L6D3_ToMinus(
.data_in(MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus),
.enable(MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus_wr_en),
.number_out(FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L1L2_L6D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L1L2_L6D3_start),
.done(FM_L1L2_L6D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus;
wire MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus_wr_en;
wire [5:0] FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L3L4_L1D3_ToMinus_MT_Layr_Minus;
wire FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L3L4_L1D3_ToMinus(
.data_in(MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus),
.enable(MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus_wr_en),
.number_out(FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L3L4_L1D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L3L4_L1D3_start),
.done(FM_L3L4_L1D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus;
wire MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus_wr_en;
wire [5:0] FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L3L4_L2D3_ToMinus_MT_Layr_Minus;
wire FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L3L4_L2D3_ToMinus(
.data_in(MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus),
.enable(MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus_wr_en),
.number_out(FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L3L4_L2D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L3L4_L2D3_start),
.done(FM_L3L4_L2D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus;
wire MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus_wr_en;
wire [5:0] FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L3L4_L5D3_ToMinus_MT_Layr_Minus;
wire FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L3L4_L5D3_ToMinus(
.data_in(MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus),
.enable(MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus_wr_en),
.number_out(FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L3L4_L5D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L3L4_L5D3_start),
.done(FM_L3L4_L5D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus;
wire MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus_wr_en;
wire [5:0] FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L3L4_L6D3_ToMinus_MT_Layr_Minus;
wire FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L3L4_L6D3_ToMinus(
.data_in(MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus),
.enable(MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus_wr_en),
.number_out(FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L3L4_L6D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L3L4_L6D3_start),
.done(FM_L3L4_L6D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus;
wire MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus_wr_en;
wire [5:0] FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L5L6_L1D3_ToMinus_MT_Layr_Minus;
wire FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L5L6_L1D3_ToMinus(
.data_in(MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus),
.enable(MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus_wr_en),
.number_out(FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L5L6_L1D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L5L6_L1D3_start),
.done(FM_L5L6_L1D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus;
wire MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus_wr_en;
wire [5:0] FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L5L6_L2D3_ToMinus_MT_Layr_Minus;
wire FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L5L6_L2D3_ToMinus(
.data_in(MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus),
.enable(MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus_wr_en),
.number_out(FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L5L6_L2D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L5L6_L2D3_start),
.done(FM_L5L6_L2D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus;
wire MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus_wr_en;
wire [5:0] FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L5L6_L3D3_ToMinus_MT_Layr_Minus;
wire FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L5L6_L3D3_ToMinus(
.data_in(MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus),
.enable(MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus_wr_en),
.number_out(FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L5L6_L3D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L5L6_L3D3_start),
.done(FM_L5L6_L3D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus;
wire MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus_wr_en;
wire [5:0] FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L5L6_L4D3_ToMinus_MT_Layr_Minus;
wire FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L5L6_L4D3_ToMinus(
.data_in(MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus),
.enable(MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus_wr_en),
.number_out(FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L5L6_L4D3_ToMinus_MT_Layr_Minus),
.read_en(FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L5L6_L4D3_start),
.done(FM_L5L6_L4D3_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus;
wire MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus_wr_en;
wire [5:0] FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L1L2_L3D4_ToMinus_MT_Layr_Minus;
wire FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L1L2_L3D4_ToMinus(
.data_in(MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus),
.enable(MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus_wr_en),
.number_out(FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L1L2_L3D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L1L2_L3D4_start),
.done(FM_L1L2_L3D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus;
wire MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus_wr_en;
wire [5:0] FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L1L2_L4D4_ToMinus_MT_Layr_Minus;
wire FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L1L2_L4D4_ToMinus(
.data_in(MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus),
.enable(MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus_wr_en),
.number_out(FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L1L2_L4D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L1L2_L4D4_start),
.done(FM_L1L2_L4D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus;
wire MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus_wr_en;
wire [5:0] FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L1L2_L5D4_ToMinus_MT_Layr_Minus;
wire FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L1L2_L5D4_ToMinus(
.data_in(MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus),
.enable(MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus_wr_en),
.number_out(FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L1L2_L5D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L1L2_L5D4_start),
.done(FM_L1L2_L5D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus;
wire MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus_wr_en;
wire [5:0] FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L1L2_L6D4_ToMinus_MT_Layr_Minus;
wire FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L1L2_L6D4_ToMinus(
.data_in(MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus),
.enable(MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus_wr_en),
.number_out(FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L1L2_L6D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L1L2_L6D4_start),
.done(FM_L1L2_L6D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus;
wire MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus_wr_en;
wire [5:0] FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L3L4_L1D4_ToMinus_MT_Layr_Minus;
wire FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L3L4_L1D4_ToMinus(
.data_in(MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus),
.enable(MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus_wr_en),
.number_out(FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L3L4_L1D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L3L4_L1D4_start),
.done(FM_L3L4_L1D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus;
wire MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus_wr_en;
wire [5:0] FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L3L4_L2D4_ToMinus_MT_Layr_Minus;
wire FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L3L4_L2D4_ToMinus(
.data_in(MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus),
.enable(MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus_wr_en),
.number_out(FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L3L4_L2D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L3L4_L2D4_start),
.done(FM_L3L4_L2D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus;
wire MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus_wr_en;
wire [5:0] FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L3L4_L5D4_ToMinus_MT_Layr_Minus;
wire FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L3L4_L5D4_ToMinus(
.data_in(MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus),
.enable(MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus_wr_en),
.number_out(FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L3L4_L5D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L3L4_L5D4_start),
.done(FM_L3L4_L5D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus;
wire MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus_wr_en;
wire [5:0] FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L3L4_L6D4_ToMinus_MT_Layr_Minus;
wire FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L3L4_L6D4_ToMinus(
.data_in(MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus),
.enable(MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus_wr_en),
.number_out(FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L3L4_L6D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L3L4_L6D4_start),
.done(FM_L3L4_L6D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus;
wire MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus_wr_en;
wire [5:0] FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L5L6_L1D4_ToMinus_MT_Layr_Minus;
wire FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L5L6_L1D4_ToMinus(
.data_in(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus),
.enable(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus_wr_en),
.number_out(FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L5L6_L1D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L5L6_L1D4_start),
.done(FM_L5L6_L1D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus;
wire MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus_wr_en;
wire [5:0] FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L5L6_L2D4_ToMinus_MT_Layr_Minus;
wire FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L5L6_L2D4_ToMinus(
.data_in(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus),
.enable(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus_wr_en),
.number_out(FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L5L6_L2D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L5L6_L2D4_start),
.done(FM_L5L6_L2D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus;
wire MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus_wr_en;
wire [5:0] FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L5L6_L3D4_ToMinus_MT_Layr_Minus;
wire FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L5L6_L3D4_ToMinus(
.data_in(MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus),
.enable(MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus_wr_en),
.number_out(FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L5L6_L3D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L5L6_L3D4_start),
.done(FM_L5L6_L3D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus;
wire MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus_wr_en;
wire [5:0] FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_number;
wire [9:0] FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_read_add;
wire [39:0] FM_L5L6_L4D4_ToMinus_MT_Layr_Minus;
wire FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_read_en;
FullMatch #(64) FM_L5L6_L4D4_ToMinus(
.data_in(MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus),
.enable(MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus_wr_en),
.number_out(FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_number),
.read_add(FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_read_add),
.data_out(FM_L5L6_L4D4_ToMinus_MT_Layr_Minus),
.read_en(FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_read_en),
.start(MC_L5L6_L4D4_start),
.done(FM_L5L6_L4D4_ToMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus;
wire MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus_wr_en;
wire [5:0] FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L1L2_L3D3_ToPlus_MT_Layr_Plus;
wire FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L1L2_L3D3_ToPlus(
.data_in(MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus),
.enable(MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus_wr_en),
.number_out(FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L1L2_L3D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L1L2_L3D3_start),
.done(FM_L1L2_L3D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus;
wire MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus_wr_en;
wire [5:0] FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L1L2_L4D3_ToPlus_MT_Layr_Plus;
wire FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L1L2_L4D3_ToPlus(
.data_in(MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus),
.enable(MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus_wr_en),
.number_out(FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L1L2_L4D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L1L2_L4D3_start),
.done(FM_L1L2_L4D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus;
wire MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus_wr_en;
wire [5:0] FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L1L2_L5D3_ToPlus_MT_Layr_Plus;
wire FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L1L2_L5D3_ToPlus(
.data_in(MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus),
.enable(MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus_wr_en),
.number_out(FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L1L2_L5D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L1L2_L5D3_start),
.done(FM_L1L2_L5D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus;
wire MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus_wr_en;
wire [5:0] FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L1L2_L6D3_ToPlus_MT_Layr_Plus;
wire FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L1L2_L6D3_ToPlus(
.data_in(MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus),
.enable(MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus_wr_en),
.number_out(FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L1L2_L6D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L1L2_L6D3_start),
.done(FM_L1L2_L6D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus;
wire MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus_wr_en;
wire [5:0] FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L3L4_L1D3_ToPlus_MT_Layr_Plus;
wire FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L3L4_L1D3_ToPlus(
.data_in(MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus),
.enable(MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus_wr_en),
.number_out(FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L3L4_L1D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L3L4_L1D3_start),
.done(FM_L3L4_L1D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus;
wire MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus_wr_en;
wire [5:0] FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L3L4_L2D3_ToPlus_MT_Layr_Plus;
wire FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L3L4_L2D3_ToPlus(
.data_in(MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus),
.enable(MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus_wr_en),
.number_out(FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L3L4_L2D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L3L4_L2D3_start),
.done(FM_L3L4_L2D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus;
wire MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus_wr_en;
wire [5:0] FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L3L4_L5D3_ToPlus_MT_Layr_Plus;
wire FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L3L4_L5D3_ToPlus(
.data_in(MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus),
.enable(MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus_wr_en),
.number_out(FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L3L4_L5D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L3L4_L5D3_start),
.done(FM_L3L4_L5D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus;
wire MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus_wr_en;
wire [5:0] FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L3L4_L6D3_ToPlus_MT_Layr_Plus;
wire FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L3L4_L6D3_ToPlus(
.data_in(MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus),
.enable(MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus_wr_en),
.number_out(FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L3L4_L6D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L3L4_L6D3_start),
.done(FM_L3L4_L6D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus;
wire MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus_wr_en;
wire [5:0] FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L5L6_L1D3_ToPlus_MT_Layr_Plus;
wire FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L5L6_L1D3_ToPlus(
.data_in(MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus),
.enable(MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus_wr_en),
.number_out(FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L5L6_L1D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L5L6_L1D3_start),
.done(FM_L5L6_L1D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus;
wire MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus_wr_en;
wire [5:0] FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L5L6_L2D3_ToPlus_MT_Layr_Plus;
wire FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L5L6_L2D3_ToPlus(
.data_in(MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus),
.enable(MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus_wr_en),
.number_out(FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L5L6_L2D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L5L6_L2D3_start),
.done(FM_L5L6_L2D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus;
wire MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus_wr_en;
wire [5:0] FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L5L6_L3D3_ToPlus_MT_Layr_Plus;
wire FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L5L6_L3D3_ToPlus(
.data_in(MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus),
.enable(MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus_wr_en),
.number_out(FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L5L6_L3D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L5L6_L3D3_start),
.done(FM_L5L6_L3D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus;
wire MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus_wr_en;
wire [5:0] FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L5L6_L4D3_ToPlus_MT_Layr_Plus;
wire FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L5L6_L4D3_ToPlus(
.data_in(MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus),
.enable(MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus_wr_en),
.number_out(FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L5L6_L4D3_ToPlus_MT_Layr_Plus),
.read_en(FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L5L6_L4D3_start),
.done(FM_L5L6_L4D3_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus;
wire MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus_wr_en;
wire [5:0] FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L1L2_L3D4_ToPlus_MT_Layr_Plus;
wire FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L1L2_L3D4_ToPlus(
.data_in(MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus),
.enable(MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus_wr_en),
.number_out(FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L1L2_L3D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L1L2_L3D4_start),
.done(FM_L1L2_L3D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus;
wire MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus_wr_en;
wire [5:0] FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L1L2_L4D4_ToPlus_MT_Layr_Plus;
wire FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L1L2_L4D4_ToPlus(
.data_in(MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus),
.enable(MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus_wr_en),
.number_out(FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L1L2_L4D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L1L2_L4D4_start),
.done(FM_L1L2_L4D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus;
wire MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus_wr_en;
wire [5:0] FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L1L2_L5D4_ToPlus_MT_Layr_Plus;
wire FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L1L2_L5D4_ToPlus(
.data_in(MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus),
.enable(MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus_wr_en),
.number_out(FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L1L2_L5D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L1L2_L5D4_start),
.done(FM_L1L2_L5D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus;
wire MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus_wr_en;
wire [5:0] FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L1L2_L6D4_ToPlus_MT_Layr_Plus;
wire FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L1L2_L6D4_ToPlus(
.data_in(MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus),
.enable(MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus_wr_en),
.number_out(FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L1L2_L6D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L1L2_L6D4_start),
.done(FM_L1L2_L6D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus;
wire MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus_wr_en;
wire [5:0] FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L3L4_L1D4_ToPlus_MT_Layr_Plus;
wire FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L3L4_L1D4_ToPlus(
.data_in(MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus),
.enable(MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus_wr_en),
.number_out(FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L3L4_L1D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L3L4_L1D4_start),
.done(FM_L3L4_L1D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus;
wire MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus_wr_en;
wire [5:0] FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L3L4_L2D4_ToPlus_MT_Layr_Plus;
wire FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L3L4_L2D4_ToPlus(
.data_in(MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus),
.enable(MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus_wr_en),
.number_out(FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L3L4_L2D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L3L4_L2D4_start),
.done(FM_L3L4_L2D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus;
wire MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus_wr_en;
wire [5:0] FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L3L4_L5D4_ToPlus_MT_Layr_Plus;
wire FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L3L4_L5D4_ToPlus(
.data_in(MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus),
.enable(MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus_wr_en),
.number_out(FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L3L4_L5D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L3L4_L5D4_start),
.done(FM_L3L4_L5D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus;
wire MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus_wr_en;
wire [5:0] FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L3L4_L6D4_ToPlus_MT_Layr_Plus;
wire FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L3L4_L6D4_ToPlus(
.data_in(MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus),
.enable(MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus_wr_en),
.number_out(FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L3L4_L6D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L3L4_L6D4_start),
.done(FM_L3L4_L6D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus;
wire MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus_wr_en;
wire [5:0] FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L5L6_L1D4_ToPlus_MT_Layr_Plus;
wire FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L5L6_L1D4_ToPlus(
.data_in(MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus),
.enable(MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus_wr_en),
.number_out(FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L5L6_L1D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L5L6_L1D4_start),
.done(FM_L5L6_L1D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus;
wire MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus_wr_en;
wire [5:0] FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L5L6_L2D4_ToPlus_MT_Layr_Plus;
wire FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L5L6_L2D4_ToPlus(
.data_in(MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus),
.enable(MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus_wr_en),
.number_out(FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L5L6_L2D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L5L6_L2D4_start),
.done(FM_L5L6_L2D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus;
wire MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus_wr_en;
wire [5:0] FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L5L6_L3D4_ToPlus_MT_Layr_Plus;
wire FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L5L6_L3D4_ToPlus(
.data_in(MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus),
.enable(MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus_wr_en),
.number_out(FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L5L6_L3D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L5L6_L3D4_start),
.done(FM_L5L6_L3D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus;
wire MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus_wr_en;
wire [5:0] FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_number;
wire [9:0] FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_read_add;
wire [39:0] FM_L5L6_L4D4_ToPlus_MT_Layr_Plus;
wire FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_read_en;
FullMatch #(64) FM_L5L6_L4D4_ToPlus(
.data_in(MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus),
.enable(MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus_wr_en),
.number_out(FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_number),
.read_add(FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_read_add),
.data_out(FM_L5L6_L4D4_ToPlus_MT_Layr_Plus),
.read_en(FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_read_en),
.start(MC_L5L6_L4D4_start),
.done(FM_L5L6_L4D4_ToPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L3D3_FM_L1L2_L3D3;
wire MC_L1L2_L3D3_FM_L1L2_L3D3_wr_en;
wire [5:0] FM_L1L2_L3D3_FT_L1L2_number;
wire [9:0] FM_L1L2_L3D3_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L3D3_FT_L1L2;
wire FM_L1L2_L3D3_FT_L1L2_read_en;
FullMatch  FM_L1L2_L3D3(
.data_in(MC_L1L2_L3D3_FM_L1L2_L3D3),
.enable(MC_L1L2_L3D3_FM_L1L2_L3D3_wr_en),
.number_out(FM_L1L2_L3D3_FT_L1L2_number),
.read_add(FM_L1L2_L3D3_FT_L1L2_read_add),
.data_out(FM_L1L2_L3D3_FT_L1L2),
.read_en(FM_L1L2_L3D3_FT_L1L2_read_en),
.start(MC_L1L2_L3D3_start),
.done(FM_L1L2_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L3D4_FM_L1L2_L3D4;
wire MC_L1L2_L3D4_FM_L1L2_L3D4_wr_en;
wire [5:0] FM_L1L2_L3D4_FT_L1L2_number;
wire [9:0] FM_L1L2_L3D4_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L3D4_FT_L1L2;
wire FM_L1L2_L3D4_FT_L1L2_read_en;
FullMatch  FM_L1L2_L3D4(
.data_in(MC_L1L2_L3D4_FM_L1L2_L3D4),
.enable(MC_L1L2_L3D4_FM_L1L2_L3D4_wr_en),
.number_out(FM_L1L2_L3D4_FT_L1L2_number),
.read_add(FM_L1L2_L3D4_FT_L1L2_read_add),
.data_out(FM_L1L2_L3D4_FT_L1L2),
.read_en(FM_L1L2_L3D4_FT_L1L2_read_en),
.start(MC_L1L2_L3D4_start),
.done(FM_L1L2_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L4D3_FM_L1L2_L4D3;
wire MC_L1L2_L4D3_FM_L1L2_L4D3_wr_en;
wire [5:0] FM_L1L2_L4D3_FT_L1L2_number;
wire [9:0] FM_L1L2_L4D3_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L4D3_FT_L1L2;
wire FM_L1L2_L4D3_FT_L1L2_read_en;
FullMatch  FM_L1L2_L4D3(
.data_in(MC_L1L2_L4D3_FM_L1L2_L4D3),
.enable(MC_L1L2_L4D3_FM_L1L2_L4D3_wr_en),
.number_out(FM_L1L2_L4D3_FT_L1L2_number),
.read_add(FM_L1L2_L4D3_FT_L1L2_read_add),
.data_out(FM_L1L2_L4D3_FT_L1L2),
.read_en(FM_L1L2_L4D3_FT_L1L2_read_en),
.start(MC_L1L2_L4D3_start),
.done(FM_L1L2_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L4D4_FM_L1L2_L4D4;
wire MC_L1L2_L4D4_FM_L1L2_L4D4_wr_en;
wire [5:0] FM_L1L2_L4D4_FT_L1L2_number;
wire [9:0] FM_L1L2_L4D4_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L4D4_FT_L1L2;
wire FM_L1L2_L4D4_FT_L1L2_read_en;
FullMatch  FM_L1L2_L4D4(
.data_in(MC_L1L2_L4D4_FM_L1L2_L4D4),
.enable(MC_L1L2_L4D4_FM_L1L2_L4D4_wr_en),
.number_out(FM_L1L2_L4D4_FT_L1L2_number),
.read_add(FM_L1L2_L4D4_FT_L1L2_read_add),
.data_out(FM_L1L2_L4D4_FT_L1L2),
.read_en(FM_L1L2_L4D4_FT_L1L2_read_en),
.start(MC_L1L2_L4D4_start),
.done(FM_L1L2_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L5D3_FM_L1L2_L5D3;
wire MC_L1L2_L5D3_FM_L1L2_L5D3_wr_en;
wire [5:0] FM_L1L2_L5D3_FT_L1L2_number;
wire [9:0] FM_L1L2_L5D3_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L5D3_FT_L1L2;
wire FM_L1L2_L5D3_FT_L1L2_read_en;
FullMatch  FM_L1L2_L5D3(
.data_in(MC_L1L2_L5D3_FM_L1L2_L5D3),
.enable(MC_L1L2_L5D3_FM_L1L2_L5D3_wr_en),
.number_out(FM_L1L2_L5D3_FT_L1L2_number),
.read_add(FM_L1L2_L5D3_FT_L1L2_read_add),
.data_out(FM_L1L2_L5D3_FT_L1L2),
.read_en(FM_L1L2_L5D3_FT_L1L2_read_en),
.start(MC_L1L2_L5D3_start),
.done(FM_L1L2_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L5D4_FM_L1L2_L5D4;
wire MC_L1L2_L5D4_FM_L1L2_L5D4_wr_en;
wire [5:0] FM_L1L2_L5D4_FT_L1L2_number;
wire [9:0] FM_L1L2_L5D4_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L5D4_FT_L1L2;
wire FM_L1L2_L5D4_FT_L1L2_read_en;
FullMatch  FM_L1L2_L5D4(
.data_in(MC_L1L2_L5D4_FM_L1L2_L5D4),
.enable(MC_L1L2_L5D4_FM_L1L2_L5D4_wr_en),
.number_out(FM_L1L2_L5D4_FT_L1L2_number),
.read_add(FM_L1L2_L5D4_FT_L1L2_read_add),
.data_out(FM_L1L2_L5D4_FT_L1L2),
.read_en(FM_L1L2_L5D4_FT_L1L2_read_en),
.start(MC_L1L2_L5D4_start),
.done(FM_L1L2_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L6D3_FM_L1L2_L6D3;
wire MC_L1L2_L6D3_FM_L1L2_L6D3_wr_en;
wire [5:0] FM_L1L2_L6D3_FT_L1L2_number;
wire [9:0] FM_L1L2_L6D3_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L6D3_FT_L1L2;
wire FM_L1L2_L6D3_FT_L1L2_read_en;
FullMatch  FM_L1L2_L6D3(
.data_in(MC_L1L2_L6D3_FM_L1L2_L6D3),
.enable(MC_L1L2_L6D3_FM_L1L2_L6D3_wr_en),
.number_out(FM_L1L2_L6D3_FT_L1L2_number),
.read_add(FM_L1L2_L6D3_FT_L1L2_read_add),
.data_out(FM_L1L2_L6D3_FT_L1L2),
.read_en(FM_L1L2_L6D3_FT_L1L2_read_en),
.start(MC_L1L2_L6D3_start),
.done(FM_L1L2_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L1L2_L6D4_FM_L1L2_L6D4;
wire MC_L1L2_L6D4_FM_L1L2_L6D4_wr_en;
wire [5:0] FM_L1L2_L6D4_FT_L1L2_number;
wire [9:0] FM_L1L2_L6D4_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L6D4_FT_L1L2;
wire FM_L1L2_L6D4_FT_L1L2_read_en;
FullMatch  FM_L1L2_L6D4(
.data_in(MC_L1L2_L6D4_FM_L1L2_L6D4),
.enable(MC_L1L2_L6D4_FM_L1L2_L6D4_wr_en),
.number_out(FM_L1L2_L6D4_FT_L1L2_number),
.read_add(FM_L1L2_L6D4_FT_L1L2_read_add),
.data_out(FM_L1L2_L6D4_FT_L1L2),
.read_en(FM_L1L2_L6D4_FT_L1L2_read_en),
.start(MC_L1L2_L6D4_start),
.done(FM_L1L2_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L1D3L2D3_TPAR_L1D3L2D3;
wire TC_L1D3L2D3_TPAR_L1D3L2D3_wr_en;
wire [10:0] TPAR_L1D3L2D3_FT_L1L2_read_add;
wire [67:0] TPAR_L1D3L2D3_FT_L1L2;
TrackletParameters  TPAR_L1D3L2D3(
.data_in(TC_L1D3L2D3_TPAR_L1D3L2D3),
.enable(TC_L1D3L2D3_TPAR_L1D3L2D3_wr_en),
.read_add(TPAR_L1D3L2D3_FT_L1L2_read_add),
.data_out(TPAR_L1D3L2D3_FT_L1L2),
.start(TC_L1D3L2D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L1D3L2D4_TPAR_L1D3L2D4;
wire TC_L1D3L2D4_TPAR_L1D3L2D4_wr_en;
wire [10:0] TPAR_L1D3L2D4_FT_L1L2_read_add;
wire [67:0] TPAR_L1D3L2D4_FT_L1L2;
TrackletParameters  TPAR_L1D3L2D4(
.data_in(TC_L1D3L2D4_TPAR_L1D3L2D4),
.enable(TC_L1D3L2D4_TPAR_L1D3L2D4_wr_en),
.read_add(TPAR_L1D3L2D4_FT_L1L2_read_add),
.data_out(TPAR_L1D3L2D4_FT_L1L2),
.start(TC_L1D3L2D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L1D4L2D4_TPAR_L1D4L2D4;
wire TC_L1D4L2D4_TPAR_L1D4L2D4_wr_en;
wire [10:0] TPAR_L1D4L2D4_FT_L1L2_read_add;
wire [67:0] TPAR_L1D4L2D4_FT_L1L2;
TrackletParameters  TPAR_L1D4L2D4(
.data_in(TC_L1D4L2D4_TPAR_L1D4L2D4),
.enable(TC_L1D4L2D4_TPAR_L1D4L2D4_wr_en),
.read_add(TPAR_L1D4L2D4_FT_L1L2_read_add),
.data_out(TPAR_L1D4L2D4_FT_L1L2),
.start(TC_L1D4L2D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L1L2_L3_FromPlus;
wire MT_Layr_Plus_FM_L1L2_L3_FromPlus_wr_en;
wire [5:0] FM_L1L2_L3_FromPlus_FT_L1L2_number;
wire [9:0] FM_L1L2_L3_FromPlus_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L3_FromPlus_FT_L1L2;
wire FM_L1L2_L3_FromPlus_FT_L1L2_read_en;
FullMatch #(64) FM_L1L2_L3_FromPlus(
.data_in(MT_Layr_Plus_FM_L1L2_L3_FromPlus),
.enable(MT_Layr_Plus_FM_L1L2_L3_FromPlus_wr_en),
.number_out(FM_L1L2_L3_FromPlus_FT_L1L2_number),
.read_add(FM_L1L2_L3_FromPlus_FT_L1L2_read_add),
.data_out(FM_L1L2_L3_FromPlus_FT_L1L2),
.read_en(FM_L1L2_L3_FromPlus_FT_L1L2_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L1L2_L3_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L1L2_L4_FromPlus;
wire MT_Layr_Plus_FM_L1L2_L4_FromPlus_wr_en;
wire [5:0] FM_L1L2_L4_FromPlus_FT_L1L2_number;
wire [9:0] FM_L1L2_L4_FromPlus_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L4_FromPlus_FT_L1L2;
wire FM_L1L2_L4_FromPlus_FT_L1L2_read_en;
FullMatch #(64) FM_L1L2_L4_FromPlus(
.data_in(MT_Layr_Plus_FM_L1L2_L4_FromPlus),
.enable(MT_Layr_Plus_FM_L1L2_L4_FromPlus_wr_en),
.number_out(FM_L1L2_L4_FromPlus_FT_L1L2_number),
.read_add(FM_L1L2_L4_FromPlus_FT_L1L2_read_add),
.data_out(FM_L1L2_L4_FromPlus_FT_L1L2),
.read_en(FM_L1L2_L4_FromPlus_FT_L1L2_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L1L2_L4_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L1L2_L5_FromPlus;
wire MT_Layr_Plus_FM_L1L2_L5_FromPlus_wr_en;
wire [5:0] FM_L1L2_L5_FromPlus_FT_L1L2_number;
wire [9:0] FM_L1L2_L5_FromPlus_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L5_FromPlus_FT_L1L2;
wire FM_L1L2_L5_FromPlus_FT_L1L2_read_en;
FullMatch #(64) FM_L1L2_L5_FromPlus(
.data_in(MT_Layr_Plus_FM_L1L2_L5_FromPlus),
.enable(MT_Layr_Plus_FM_L1L2_L5_FromPlus_wr_en),
.number_out(FM_L1L2_L5_FromPlus_FT_L1L2_number),
.read_add(FM_L1L2_L5_FromPlus_FT_L1L2_read_add),
.data_out(FM_L1L2_L5_FromPlus_FT_L1L2),
.read_en(FM_L1L2_L5_FromPlus_FT_L1L2_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L1L2_L5_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L1L2_L6_FromPlus;
wire MT_Layr_Plus_FM_L1L2_L6_FromPlus_wr_en;
wire [5:0] FM_L1L2_L6_FromPlus_FT_L1L2_number;
wire [9:0] FM_L1L2_L6_FromPlus_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L6_FromPlus_FT_L1L2;
wire FM_L1L2_L6_FromPlus_FT_L1L2_read_en;
FullMatch #(64) FM_L1L2_L6_FromPlus(
.data_in(MT_Layr_Plus_FM_L1L2_L6_FromPlus),
.enable(MT_Layr_Plus_FM_L1L2_L6_FromPlus_wr_en),
.number_out(FM_L1L2_L6_FromPlus_FT_L1L2_number),
.read_add(FM_L1L2_L6_FromPlus_FT_L1L2_read_add),
.data_out(FM_L1L2_L6_FromPlus_FT_L1L2),
.read_en(FM_L1L2_L6_FromPlus_FT_L1L2_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L1L2_L6_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L1L2_L3_FromMinus;
wire MT_Layr_Minus_FM_L1L2_L3_FromMinus_wr_en;
wire [5:0] FM_L1L2_L3_FromMinus_FT_L1L2_number;
wire [9:0] FM_L1L2_L3_FromMinus_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L3_FromMinus_FT_L1L2;
wire FM_L1L2_L3_FromMinus_FT_L1L2_read_en;
FullMatch #(64) FM_L1L2_L3_FromMinus(
.data_in(MT_Layr_Minus_FM_L1L2_L3_FromMinus),
.enable(MT_Layr_Minus_FM_L1L2_L3_FromMinus_wr_en),
.number_out(FM_L1L2_L3_FromMinus_FT_L1L2_number),
.read_add(FM_L1L2_L3_FromMinus_FT_L1L2_read_add),
.data_out(FM_L1L2_L3_FromMinus_FT_L1L2),
.read_en(FM_L1L2_L3_FromMinus_FT_L1L2_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L1L2_L3_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L1L2_L4_FromMinus;
wire MT_Layr_Minus_FM_L1L2_L4_FromMinus_wr_en;
wire [5:0] FM_L1L2_L4_FromMinus_FT_L1L2_number;
wire [9:0] FM_L1L2_L4_FromMinus_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L4_FromMinus_FT_L1L2;
wire FM_L1L2_L4_FromMinus_FT_L1L2_read_en;
FullMatch #(64) FM_L1L2_L4_FromMinus(
.data_in(MT_Layr_Minus_FM_L1L2_L4_FromMinus),
.enable(MT_Layr_Minus_FM_L1L2_L4_FromMinus_wr_en),
.number_out(FM_L1L2_L4_FromMinus_FT_L1L2_number),
.read_add(FM_L1L2_L4_FromMinus_FT_L1L2_read_add),
.data_out(FM_L1L2_L4_FromMinus_FT_L1L2),
.read_en(FM_L1L2_L4_FromMinus_FT_L1L2_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L1L2_L4_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L1L2_L5_FromMinus;
wire MT_Layr_Minus_FM_L1L2_L5_FromMinus_wr_en;
wire [5:0] FM_L1L2_L5_FromMinus_FT_L1L2_number;
wire [9:0] FM_L1L2_L5_FromMinus_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L5_FromMinus_FT_L1L2;
wire FM_L1L2_L5_FromMinus_FT_L1L2_read_en;
FullMatch #(64) FM_L1L2_L5_FromMinus(
.data_in(MT_Layr_Minus_FM_L1L2_L5_FromMinus),
.enable(MT_Layr_Minus_FM_L1L2_L5_FromMinus_wr_en),
.number_out(FM_L1L2_L5_FromMinus_FT_L1L2_number),
.read_add(FM_L1L2_L5_FromMinus_FT_L1L2_read_add),
.data_out(FM_L1L2_L5_FromMinus_FT_L1L2),
.read_en(FM_L1L2_L5_FromMinus_FT_L1L2_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L1L2_L5_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L1L2_L6_FromMinus;
wire MT_Layr_Minus_FM_L1L2_L6_FromMinus_wr_en;
wire [5:0] FM_L1L2_L6_FromMinus_FT_L1L2_number;
wire [9:0] FM_L1L2_L6_FromMinus_FT_L1L2_read_add;
wire [39:0] FM_L1L2_L6_FromMinus_FT_L1L2;
wire FM_L1L2_L6_FromMinus_FT_L1L2_read_en;
FullMatch #(64) FM_L1L2_L6_FromMinus(
.data_in(MT_Layr_Minus_FM_L1L2_L6_FromMinus),
.enable(MT_Layr_Minus_FM_L1L2_L6_FromMinus_wr_en),
.number_out(FM_L1L2_L6_FromMinus_FT_L1L2_number),
.read_add(FM_L1L2_L6_FromMinus_FT_L1L2_read_add),
.data_out(FM_L1L2_L6_FromMinus_FT_L1L2),
.read_en(FM_L1L2_L6_FromMinus_FT_L1L2_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L1L2_L6_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L1D3_FM_L3L4_L1D3;
wire MC_L3L4_L1D3_FM_L3L4_L1D3_wr_en;
wire [5:0] FM_L3L4_L1D3_FT_L3L4_number;
wire [9:0] FM_L3L4_L1D3_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L1D3_FT_L3L4;
wire FM_L3L4_L1D3_FT_L3L4_read_en;
FullMatch  FM_L3L4_L1D3(
.data_in(MC_L3L4_L1D3_FM_L3L4_L1D3),
.enable(MC_L3L4_L1D3_FM_L3L4_L1D3_wr_en),
.number_out(FM_L3L4_L1D3_FT_L3L4_number),
.read_add(FM_L3L4_L1D3_FT_L3L4_read_add),
.data_out(FM_L3L4_L1D3_FT_L3L4),
.read_en(FM_L3L4_L1D3_FT_L3L4_read_en),
.start(MC_L3L4_L1D3_start),
.done(FM_L3L4_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L1D4_FM_L3L4_L1D4;
wire MC_L3L4_L1D4_FM_L3L4_L1D4_wr_en;
wire [5:0] FM_L3L4_L1D4_FT_L3L4_number;
wire [9:0] FM_L3L4_L1D4_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L1D4_FT_L3L4;
wire FM_L3L4_L1D4_FT_L3L4_read_en;
FullMatch  FM_L3L4_L1D4(
.data_in(MC_L3L4_L1D4_FM_L3L4_L1D4),
.enable(MC_L3L4_L1D4_FM_L3L4_L1D4_wr_en),
.number_out(FM_L3L4_L1D4_FT_L3L4_number),
.read_add(FM_L3L4_L1D4_FT_L3L4_read_add),
.data_out(FM_L3L4_L1D4_FT_L3L4),
.read_en(FM_L3L4_L1D4_FT_L3L4_read_en),
.start(MC_L3L4_L1D4_start),
.done(FM_L3L4_L1D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L2D3_FM_L3L4_L2D3;
wire MC_L3L4_L2D3_FM_L3L4_L2D3_wr_en;
wire [5:0] FM_L3L4_L2D3_FT_L3L4_number;
wire [9:0] FM_L3L4_L2D3_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L2D3_FT_L3L4;
wire FM_L3L4_L2D3_FT_L3L4_read_en;
FullMatch  FM_L3L4_L2D3(
.data_in(MC_L3L4_L2D3_FM_L3L4_L2D3),
.enable(MC_L3L4_L2D3_FM_L3L4_L2D3_wr_en),
.number_out(FM_L3L4_L2D3_FT_L3L4_number),
.read_add(FM_L3L4_L2D3_FT_L3L4_read_add),
.data_out(FM_L3L4_L2D3_FT_L3L4),
.read_en(FM_L3L4_L2D3_FT_L3L4_read_en),
.start(MC_L3L4_L2D3_start),
.done(FM_L3L4_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L2D4_FM_L3L4_L2D4;
wire MC_L3L4_L2D4_FM_L3L4_L2D4_wr_en;
wire [5:0] FM_L3L4_L2D4_FT_L3L4_number;
wire [9:0] FM_L3L4_L2D4_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L2D4_FT_L3L4;
wire FM_L3L4_L2D4_FT_L3L4_read_en;
FullMatch  FM_L3L4_L2D4(
.data_in(MC_L3L4_L2D4_FM_L3L4_L2D4),
.enable(MC_L3L4_L2D4_FM_L3L4_L2D4_wr_en),
.number_out(FM_L3L4_L2D4_FT_L3L4_number),
.read_add(FM_L3L4_L2D4_FT_L3L4_read_add),
.data_out(FM_L3L4_L2D4_FT_L3L4),
.read_en(FM_L3L4_L2D4_FT_L3L4_read_en),
.start(MC_L3L4_L2D4_start),
.done(FM_L3L4_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L5D3_FM_L3L4_L5D3;
wire MC_L3L4_L5D3_FM_L3L4_L5D3_wr_en;
wire [5:0] FM_L3L4_L5D3_FT_L3L4_number;
wire [9:0] FM_L3L4_L5D3_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L5D3_FT_L3L4;
wire FM_L3L4_L5D3_FT_L3L4_read_en;
FullMatch  FM_L3L4_L5D3(
.data_in(MC_L3L4_L5D3_FM_L3L4_L5D3),
.enable(MC_L3L4_L5D3_FM_L3L4_L5D3_wr_en),
.number_out(FM_L3L4_L5D3_FT_L3L4_number),
.read_add(FM_L3L4_L5D3_FT_L3L4_read_add),
.data_out(FM_L3L4_L5D3_FT_L3L4),
.read_en(FM_L3L4_L5D3_FT_L3L4_read_en),
.start(MC_L3L4_L5D3_start),
.done(FM_L3L4_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L5D4_FM_L3L4_L5D4;
wire MC_L3L4_L5D4_FM_L3L4_L5D4_wr_en;
wire [5:0] FM_L3L4_L5D4_FT_L3L4_number;
wire [9:0] FM_L3L4_L5D4_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L5D4_FT_L3L4;
wire FM_L3L4_L5D4_FT_L3L4_read_en;
FullMatch  FM_L3L4_L5D4(
.data_in(MC_L3L4_L5D4_FM_L3L4_L5D4),
.enable(MC_L3L4_L5D4_FM_L3L4_L5D4_wr_en),
.number_out(FM_L3L4_L5D4_FT_L3L4_number),
.read_add(FM_L3L4_L5D4_FT_L3L4_read_add),
.data_out(FM_L3L4_L5D4_FT_L3L4),
.read_en(FM_L3L4_L5D4_FT_L3L4_read_en),
.start(MC_L3L4_L5D4_start),
.done(FM_L3L4_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L6D3_FM_L3L4_L6D3;
wire MC_L3L4_L6D3_FM_L3L4_L6D3_wr_en;
wire [5:0] FM_L3L4_L6D3_FT_L3L4_number;
wire [9:0] FM_L3L4_L6D3_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L6D3_FT_L3L4;
wire FM_L3L4_L6D3_FT_L3L4_read_en;
FullMatch  FM_L3L4_L6D3(
.data_in(MC_L3L4_L6D3_FM_L3L4_L6D3),
.enable(MC_L3L4_L6D3_FM_L3L4_L6D3_wr_en),
.number_out(FM_L3L4_L6D3_FT_L3L4_number),
.read_add(FM_L3L4_L6D3_FT_L3L4_read_add),
.data_out(FM_L3L4_L6D3_FT_L3L4),
.read_en(FM_L3L4_L6D3_FT_L3L4_read_en),
.start(MC_L3L4_L6D3_start),
.done(FM_L3L4_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L3L4_L6D4_FM_L3L4_L6D4;
wire MC_L3L4_L6D4_FM_L3L4_L6D4_wr_en;
wire [5:0] FM_L3L4_L6D4_FT_L3L4_number;
wire [9:0] FM_L3L4_L6D4_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L6D4_FT_L3L4;
wire FM_L3L4_L6D4_FT_L3L4_read_en;
FullMatch  FM_L3L4_L6D4(
.data_in(MC_L3L4_L6D4_FM_L3L4_L6D4),
.enable(MC_L3L4_L6D4_FM_L3L4_L6D4_wr_en),
.number_out(FM_L3L4_L6D4_FT_L3L4_number),
.read_add(FM_L3L4_L6D4_FT_L3L4_read_add),
.data_out(FM_L3L4_L6D4_FT_L3L4),
.read_en(FM_L3L4_L6D4_FT_L3L4_read_en),
.start(MC_L3L4_L6D4_start),
.done(FM_L3L4_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L3L4_L1_FromMinus;
wire MT_Layr_Minus_FM_L3L4_L1_FromMinus_wr_en;
wire [5:0] FM_L3L4_L1_FromMinus_FT_L3L4_number;
wire [9:0] FM_L3L4_L1_FromMinus_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L1_FromMinus_FT_L3L4;
wire FM_L3L4_L1_FromMinus_FT_L3L4_read_en;
FullMatch #(64) FM_L3L4_L1_FromMinus(
.data_in(MT_Layr_Minus_FM_L3L4_L1_FromMinus),
.enable(MT_Layr_Minus_FM_L3L4_L1_FromMinus_wr_en),
.number_out(FM_L3L4_L1_FromMinus_FT_L3L4_number),
.read_add(FM_L3L4_L1_FromMinus_FT_L3L4_read_add),
.data_out(FM_L3L4_L1_FromMinus_FT_L3L4),
.read_en(FM_L3L4_L1_FromMinus_FT_L3L4_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L3L4_L1_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L3L4_L2_FromMinus;
wire MT_Layr_Minus_FM_L3L4_L2_FromMinus_wr_en;
wire [5:0] FM_L3L4_L2_FromMinus_FT_L3L4_number;
wire [9:0] FM_L3L4_L2_FromMinus_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L2_FromMinus_FT_L3L4;
wire FM_L3L4_L2_FromMinus_FT_L3L4_read_en;
FullMatch #(64) FM_L3L4_L2_FromMinus(
.data_in(MT_Layr_Minus_FM_L3L4_L2_FromMinus),
.enable(MT_Layr_Minus_FM_L3L4_L2_FromMinus_wr_en),
.number_out(FM_L3L4_L2_FromMinus_FT_L3L4_number),
.read_add(FM_L3L4_L2_FromMinus_FT_L3L4_read_add),
.data_out(FM_L3L4_L2_FromMinus_FT_L3L4),
.read_en(FM_L3L4_L2_FromMinus_FT_L3L4_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L3L4_L2_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L3L4_L5_FromMinus;
wire MT_Layr_Minus_FM_L3L4_L5_FromMinus_wr_en;
wire [5:0] FM_L3L4_L5_FromMinus_FT_L3L4_number;
wire [9:0] FM_L3L4_L5_FromMinus_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L5_FromMinus_FT_L3L4;
wire FM_L3L4_L5_FromMinus_FT_L3L4_read_en;
FullMatch #(64) FM_L3L4_L5_FromMinus(
.data_in(MT_Layr_Minus_FM_L3L4_L5_FromMinus),
.enable(MT_Layr_Minus_FM_L3L4_L5_FromMinus_wr_en),
.number_out(FM_L3L4_L5_FromMinus_FT_L3L4_number),
.read_add(FM_L3L4_L5_FromMinus_FT_L3L4_read_add),
.data_out(FM_L3L4_L5_FromMinus_FT_L3L4),
.read_en(FM_L3L4_L5_FromMinus_FT_L3L4_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L3L4_L5_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L3L4_L6_FromMinus;
wire MT_Layr_Minus_FM_L3L4_L6_FromMinus_wr_en;
wire [5:0] FM_L3L4_L6_FromMinus_FT_L3L4_number;
wire [9:0] FM_L3L4_L6_FromMinus_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L6_FromMinus_FT_L3L4;
wire FM_L3L4_L6_FromMinus_FT_L3L4_read_en;
FullMatch #(64) FM_L3L4_L6_FromMinus(
.data_in(MT_Layr_Minus_FM_L3L4_L6_FromMinus),
.enable(MT_Layr_Minus_FM_L3L4_L6_FromMinus_wr_en),
.number_out(FM_L3L4_L6_FromMinus_FT_L3L4_number),
.read_add(FM_L3L4_L6_FromMinus_FT_L3L4_read_add),
.data_out(FM_L3L4_L6_FromMinus_FT_L3L4),
.read_en(FM_L3L4_L6_FromMinus_FT_L3L4_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L3L4_L6_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L3L4_L1_FromPlus;
wire MT_Layr_Plus_FM_L3L4_L1_FromPlus_wr_en;
wire [5:0] FM_L3L4_L1_FromPlus_FT_L3L4_number;
wire [9:0] FM_L3L4_L1_FromPlus_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L1_FromPlus_FT_L3L4;
wire FM_L3L4_L1_FromPlus_FT_L3L4_read_en;
FullMatch #(64) FM_L3L4_L1_FromPlus(
.data_in(MT_Layr_Plus_FM_L3L4_L1_FromPlus),
.enable(MT_Layr_Plus_FM_L3L4_L1_FromPlus_wr_en),
.number_out(FM_L3L4_L1_FromPlus_FT_L3L4_number),
.read_add(FM_L3L4_L1_FromPlus_FT_L3L4_read_add),
.data_out(FM_L3L4_L1_FromPlus_FT_L3L4),
.read_en(FM_L3L4_L1_FromPlus_FT_L3L4_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L3L4_L1_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L3L4_L2_FromPlus;
wire MT_Layr_Plus_FM_L3L4_L2_FromPlus_wr_en;
wire [5:0] FM_L3L4_L2_FromPlus_FT_L3L4_number;
wire [9:0] FM_L3L4_L2_FromPlus_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L2_FromPlus_FT_L3L4;
wire FM_L3L4_L2_FromPlus_FT_L3L4_read_en;
FullMatch #(64) FM_L3L4_L2_FromPlus(
.data_in(MT_Layr_Plus_FM_L3L4_L2_FromPlus),
.enable(MT_Layr_Plus_FM_L3L4_L2_FromPlus_wr_en),
.number_out(FM_L3L4_L2_FromPlus_FT_L3L4_number),
.read_add(FM_L3L4_L2_FromPlus_FT_L3L4_read_add),
.data_out(FM_L3L4_L2_FromPlus_FT_L3L4),
.read_en(FM_L3L4_L2_FromPlus_FT_L3L4_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L3L4_L2_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L3L4_L5_FromPlus;
wire MT_Layr_Plus_FM_L3L4_L5_FromPlus_wr_en;
wire [5:0] FM_L3L4_L5_FromPlus_FT_L3L4_number;
wire [9:0] FM_L3L4_L5_FromPlus_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L5_FromPlus_FT_L3L4;
wire FM_L3L4_L5_FromPlus_FT_L3L4_read_en;
FullMatch #(64) FM_L3L4_L5_FromPlus(
.data_in(MT_Layr_Plus_FM_L3L4_L5_FromPlus),
.enable(MT_Layr_Plus_FM_L3L4_L5_FromPlus_wr_en),
.number_out(FM_L3L4_L5_FromPlus_FT_L3L4_number),
.read_add(FM_L3L4_L5_FromPlus_FT_L3L4_read_add),
.data_out(FM_L3L4_L5_FromPlus_FT_L3L4),
.read_en(FM_L3L4_L5_FromPlus_FT_L3L4_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L3L4_L5_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L3L4_L6_FromPlus;
wire MT_Layr_Plus_FM_L3L4_L6_FromPlus_wr_en;
wire [5:0] FM_L3L4_L6_FromPlus_FT_L3L4_number;
wire [9:0] FM_L3L4_L6_FromPlus_FT_L3L4_read_add;
wire [39:0] FM_L3L4_L6_FromPlus_FT_L3L4;
wire FM_L3L4_L6_FromPlus_FT_L3L4_read_en;
FullMatch #(64) FM_L3L4_L6_FromPlus(
.data_in(MT_Layr_Plus_FM_L3L4_L6_FromPlus),
.enable(MT_Layr_Plus_FM_L3L4_L6_FromPlus_wr_en),
.number_out(FM_L3L4_L6_FromPlus_FT_L3L4_number),
.read_add(FM_L3L4_L6_FromPlus_FT_L3L4_read_add),
.data_out(FM_L3L4_L6_FromPlus_FT_L3L4),
.read_en(FM_L3L4_L6_FromPlus_FT_L3L4_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L3L4_L6_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L3D3L4D3_TPAR_L3D3L4D3;
wire TC_L3D3L4D3_TPAR_L3D3L4D3_wr_en;
wire [10:0] TPAR_L3D3L4D3_FT_L3L4_read_add;
wire [67:0] TPAR_L3D3L4D3_FT_L3L4;
TrackletParameters  TPAR_L3D3L4D3(
.data_in(TC_L3D3L4D3_TPAR_L3D3L4D3),
.enable(TC_L3D3L4D3_TPAR_L3D3L4D3_wr_en),
.read_add(TPAR_L3D3L4D3_FT_L3L4_read_add),
.data_out(TPAR_L3D3L4D3_FT_L3L4),
.start(TC_L3D3L4D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L3D3L4D4_TPAR_L3D3L4D4;
wire TC_L3D3L4D4_TPAR_L3D3L4D4_wr_en;
wire [10:0] TPAR_L3D3L4D4_FT_L3L4_read_add;
wire [67:0] TPAR_L3D3L4D4_FT_L3L4;
TrackletParameters  TPAR_L3D3L4D4(
.data_in(TC_L3D3L4D4_TPAR_L3D3L4D4),
.enable(TC_L3D3L4D4_TPAR_L3D3L4D4_wr_en),
.read_add(TPAR_L3D3L4D4_FT_L3L4_read_add),
.data_out(TPAR_L3D3L4D4_FT_L3L4),
.start(TC_L3D3L4D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L3D4L4D4_TPAR_L3D4L4D4;
wire TC_L3D4L4D4_TPAR_L3D4L4D4_wr_en;
wire [10:0] TPAR_L3D4L4D4_FT_L3L4_read_add;
wire [67:0] TPAR_L3D4L4D4_FT_L3L4;
TrackletParameters  TPAR_L3D4L4D4(
.data_in(TC_L3D4L4D4_TPAR_L3D4L4D4),
.enable(TC_L3D4L4D4_TPAR_L3D4L4D4_wr_en),
.read_add(TPAR_L3D4L4D4_FT_L3L4_read_add),
.data_out(TPAR_L3D4L4D4_FT_L3L4),
.start(TC_L3D4L4D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L1D3_FM_L5L6_L1D3;
wire MC_L5L6_L1D3_FM_L5L6_L1D3_wr_en;
wire [5:0] FM_L5L6_L1D3_FT_L5L6_number;
wire [9:0] FM_L5L6_L1D3_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L1D3_FT_L5L6;
wire FM_L5L6_L1D3_FT_L5L6_read_en;
FullMatch  FM_L5L6_L1D3(
.data_in(MC_L5L6_L1D3_FM_L5L6_L1D3),
.enable(MC_L5L6_L1D3_FM_L5L6_L1D3_wr_en),
.number_out(FM_L5L6_L1D3_FT_L5L6_number),
.read_add(FM_L5L6_L1D3_FT_L5L6_read_add),
.data_out(FM_L5L6_L1D3_FT_L5L6),
.read_en(FM_L5L6_L1D3_FT_L5L6_read_en),
.start(MC_L5L6_L1D3_start),
.done(FM_L5L6_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L1D4_FM_L5L6_L1D4;
wire MC_L5L6_L1D4_FM_L5L6_L1D4_wr_en;
wire [5:0] FM_L5L6_L1D4_FT_L5L6_number;
wire [9:0] FM_L5L6_L1D4_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L1D4_FT_L5L6;
wire FM_L5L6_L1D4_FT_L5L6_read_en;
FullMatch  FM_L5L6_L1D4(
.data_in(MC_L5L6_L1D4_FM_L5L6_L1D4),
.enable(MC_L5L6_L1D4_FM_L5L6_L1D4_wr_en),
.number_out(FM_L5L6_L1D4_FT_L5L6_number),
.read_add(FM_L5L6_L1D4_FT_L5L6_read_add),
.data_out(FM_L5L6_L1D4_FT_L5L6),
.read_en(FM_L5L6_L1D4_FT_L5L6_read_en),
.start(MC_L5L6_L1D4_start),
.done(FM_L5L6_L1D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L2D3_FM_L5L6_L2D3;
wire MC_L5L6_L2D3_FM_L5L6_L2D3_wr_en;
wire [5:0] FM_L5L6_L2D3_FT_L5L6_number;
wire [9:0] FM_L5L6_L2D3_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L2D3_FT_L5L6;
wire FM_L5L6_L2D3_FT_L5L6_read_en;
FullMatch  FM_L5L6_L2D3(
.data_in(MC_L5L6_L2D3_FM_L5L6_L2D3),
.enable(MC_L5L6_L2D3_FM_L5L6_L2D3_wr_en),
.number_out(FM_L5L6_L2D3_FT_L5L6_number),
.read_add(FM_L5L6_L2D3_FT_L5L6_read_add),
.data_out(FM_L5L6_L2D3_FT_L5L6),
.read_en(FM_L5L6_L2D3_FT_L5L6_read_en),
.start(MC_L5L6_L2D3_start),
.done(FM_L5L6_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L2D4_FM_L5L6_L2D4;
wire MC_L5L6_L2D4_FM_L5L6_L2D4_wr_en;
wire [5:0] FM_L5L6_L2D4_FT_L5L6_number;
wire [9:0] FM_L5L6_L2D4_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L2D4_FT_L5L6;
wire FM_L5L6_L2D4_FT_L5L6_read_en;
FullMatch  FM_L5L6_L2D4(
.data_in(MC_L5L6_L2D4_FM_L5L6_L2D4),
.enable(MC_L5L6_L2D4_FM_L5L6_L2D4_wr_en),
.number_out(FM_L5L6_L2D4_FT_L5L6_number),
.read_add(FM_L5L6_L2D4_FT_L5L6_read_add),
.data_out(FM_L5L6_L2D4_FT_L5L6),
.read_en(FM_L5L6_L2D4_FT_L5L6_read_en),
.start(MC_L5L6_L2D4_start),
.done(FM_L5L6_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L3D3_FM_L5L6_L3D3;
wire MC_L5L6_L3D3_FM_L5L6_L3D3_wr_en;
wire [5:0] FM_L5L6_L3D3_FT_L5L6_number;
wire [9:0] FM_L5L6_L3D3_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L3D3_FT_L5L6;
wire FM_L5L6_L3D3_FT_L5L6_read_en;
FullMatch  FM_L5L6_L3D3(
.data_in(MC_L5L6_L3D3_FM_L5L6_L3D3),
.enable(MC_L5L6_L3D3_FM_L5L6_L3D3_wr_en),
.number_out(FM_L5L6_L3D3_FT_L5L6_number),
.read_add(FM_L5L6_L3D3_FT_L5L6_read_add),
.data_out(FM_L5L6_L3D3_FT_L5L6),
.read_en(FM_L5L6_L3D3_FT_L5L6_read_en),
.start(MC_L5L6_L3D3_start),
.done(FM_L5L6_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L3D4_FM_L5L6_L3D4;
wire MC_L5L6_L3D4_FM_L5L6_L3D4_wr_en;
wire [5:0] FM_L5L6_L3D4_FT_L5L6_number;
wire [9:0] FM_L5L6_L3D4_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L3D4_FT_L5L6;
wire FM_L5L6_L3D4_FT_L5L6_read_en;
FullMatch  FM_L5L6_L3D4(
.data_in(MC_L5L6_L3D4_FM_L5L6_L3D4),
.enable(MC_L5L6_L3D4_FM_L5L6_L3D4_wr_en),
.number_out(FM_L5L6_L3D4_FT_L5L6_number),
.read_add(FM_L5L6_L3D4_FT_L5L6_read_add),
.data_out(FM_L5L6_L3D4_FT_L5L6),
.read_en(FM_L5L6_L3D4_FT_L5L6_read_en),
.start(MC_L5L6_L3D4_start),
.done(FM_L5L6_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L4D3_FM_L5L6_L4D3;
wire MC_L5L6_L4D3_FM_L5L6_L4D3_wr_en;
wire [5:0] FM_L5L6_L4D3_FT_L5L6_number;
wire [9:0] FM_L5L6_L4D3_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L4D3_FT_L5L6;
wire FM_L5L6_L4D3_FT_L5L6_read_en;
FullMatch  FM_L5L6_L4D3(
.data_in(MC_L5L6_L4D3_FM_L5L6_L4D3),
.enable(MC_L5L6_L4D3_FM_L5L6_L4D3_wr_en),
.number_out(FM_L5L6_L4D3_FT_L5L6_number),
.read_add(FM_L5L6_L4D3_FT_L5L6_read_add),
.data_out(FM_L5L6_L4D3_FT_L5L6),
.read_en(FM_L5L6_L4D3_FT_L5L6_read_en),
.start(MC_L5L6_L4D3_start),
.done(FM_L5L6_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MC_L5L6_L4D4_FM_L5L6_L4D4;
wire MC_L5L6_L4D4_FM_L5L6_L4D4_wr_en;
wire [5:0] FM_L5L6_L4D4_FT_L5L6_number;
wire [9:0] FM_L5L6_L4D4_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L4D4_FT_L5L6;
wire FM_L5L6_L4D4_FT_L5L6_read_en;
FullMatch  FM_L5L6_L4D4(
.data_in(MC_L5L6_L4D4_FM_L5L6_L4D4),
.enable(MC_L5L6_L4D4_FM_L5L6_L4D4_wr_en),
.number_out(FM_L5L6_L4D4_FT_L5L6_number),
.read_add(FM_L5L6_L4D4_FT_L5L6_read_add),
.data_out(FM_L5L6_L4D4_FT_L5L6),
.read_en(FM_L5L6_L4D4_FT_L5L6_read_en),
.start(MC_L5L6_L4D4_start),
.done(FM_L5L6_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L5D3L6D3_TPAR_L5D3L6D3;
wire TC_L5D3L6D3_TPAR_L5D3L6D3_wr_en;
wire [10:0] TPAR_L5D3L6D3_FT_L5L6_read_add;
wire [67:0] TPAR_L5D3L6D3_FT_L5L6;
TrackletParameters  TPAR_L5D3L6D3(
.data_in(TC_L5D3L6D3_TPAR_L5D3L6D3),
.enable(TC_L5D3L6D3_TPAR_L5D3L6D3_wr_en),
.read_add(TPAR_L5D3L6D3_FT_L5L6_read_add),
.data_out(TPAR_L5D3L6D3_FT_L5L6),
.start(TC_L5D3L6D3_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L5D3L6D4_TPAR_L5D3L6D4;
wire TC_L5D3L6D4_TPAR_L5D3L6D4_wr_en;
wire [10:0] TPAR_L5D3L6D4_FT_L5L6_read_add;
wire [67:0] TPAR_L5D3L6D4_FT_L5L6;
TrackletParameters  TPAR_L5D3L6D4(
.data_in(TC_L5D3L6D4_TPAR_L5D3L6D4),
.enable(TC_L5D3L6D4_TPAR_L5D3L6D4_wr_en),
.read_add(TPAR_L5D3L6D4_FT_L5L6_read_add),
.data_out(TPAR_L5D3L6D4_FT_L5L6),
.start(TC_L5D3L6D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [67:0] TC_L5D4L6D4_TPAR_L5D4L6D4;
wire TC_L5D4L6D4_TPAR_L5D4L6D4_wr_en;
wire [10:0] TPAR_L5D4L6D4_FT_L5L6_read_add;
wire [67:0] TPAR_L5D4L6D4_FT_L5L6;
TrackletParameters  TPAR_L5D4L6D4(
.data_in(TC_L5D4L6D4_TPAR_L5D4L6D4),
.enable(TC_L5D4L6D4_TPAR_L5D4L6D4_wr_en),
.read_add(TPAR_L5D4L6D4_FT_L5L6_read_add),
.data_out(TPAR_L5D4L6D4_FT_L5L6),
.start(TC_L5D4L6D4_start),
.done(),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L5L6_L1_FromPlus;
wire MT_Layr_Plus_FM_L5L6_L1_FromPlus_wr_en;
wire [5:0] FM_L5L6_L1_FromPlus_FT_L5L6_number;
wire [9:0] FM_L5L6_L1_FromPlus_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L1_FromPlus_FT_L5L6;
wire FM_L5L6_L1_FromPlus_FT_L5L6_read_en;
FullMatch #(64) FM_L5L6_L1_FromPlus(
.data_in(MT_Layr_Plus_FM_L5L6_L1_FromPlus),
.enable(MT_Layr_Plus_FM_L5L6_L1_FromPlus_wr_en),
.number_out(FM_L5L6_L1_FromPlus_FT_L5L6_number),
.read_add(FM_L5L6_L1_FromPlus_FT_L5L6_read_add),
.data_out(FM_L5L6_L1_FromPlus_FT_L5L6),
.read_en(FM_L5L6_L1_FromPlus_FT_L5L6_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L5L6_L1_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L5L6_L2_FromPlus;
wire MT_Layr_Plus_FM_L5L6_L2_FromPlus_wr_en;
wire [5:0] FM_L5L6_L2_FromPlus_FT_L5L6_number;
wire [9:0] FM_L5L6_L2_FromPlus_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L2_FromPlus_FT_L5L6;
wire FM_L5L6_L2_FromPlus_FT_L5L6_read_en;
FullMatch #(64) FM_L5L6_L2_FromPlus(
.data_in(MT_Layr_Plus_FM_L5L6_L2_FromPlus),
.enable(MT_Layr_Plus_FM_L5L6_L2_FromPlus_wr_en),
.number_out(FM_L5L6_L2_FromPlus_FT_L5L6_number),
.read_add(FM_L5L6_L2_FromPlus_FT_L5L6_read_add),
.data_out(FM_L5L6_L2_FromPlus_FT_L5L6),
.read_en(FM_L5L6_L2_FromPlus_FT_L5L6_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L5L6_L2_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L5L6_L3_FromPlus;
wire MT_Layr_Plus_FM_L5L6_L3_FromPlus_wr_en;
wire [5:0] FM_L5L6_L3_FromPlus_FT_L5L6_number;
wire [9:0] FM_L5L6_L3_FromPlus_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L3_FromPlus_FT_L5L6;
wire FM_L5L6_L3_FromPlus_FT_L5L6_read_en;
FullMatch #(64) FM_L5L6_L3_FromPlus(
.data_in(MT_Layr_Plus_FM_L5L6_L3_FromPlus),
.enable(MT_Layr_Plus_FM_L5L6_L3_FromPlus_wr_en),
.number_out(FM_L5L6_L3_FromPlus_FT_L5L6_number),
.read_add(FM_L5L6_L3_FromPlus_FT_L5L6_read_add),
.data_out(FM_L5L6_L3_FromPlus_FT_L5L6),
.read_en(FM_L5L6_L3_FromPlus_FT_L5L6_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L5L6_L3_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Plus_FM_L5L6_L4_FromPlus;
wire MT_Layr_Plus_FM_L5L6_L4_FromPlus_wr_en;
wire [5:0] FM_L5L6_L4_FromPlus_FT_L5L6_number;
wire [9:0] FM_L5L6_L4_FromPlus_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L4_FromPlus_FT_L5L6;
wire FM_L5L6_L4_FromPlus_FT_L5L6_read_en;
FullMatch #(64) FM_L5L6_L4_FromPlus(
.data_in(MT_Layr_Plus_FM_L5L6_L4_FromPlus),
.enable(MT_Layr_Plus_FM_L5L6_L4_FromPlus_wr_en),
.number_out(FM_L5L6_L4_FromPlus_FT_L5L6_number),
.read_add(FM_L5L6_L4_FromPlus_FT_L5L6_read_add),
.data_out(FM_L5L6_L4_FromPlus_FT_L5L6),
.read_en(FM_L5L6_L4_FromPlus_FT_L5L6_read_en),
.start(MT_Layr_Plus_start),
.done(FM_L5L6_L4_FromPlus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L5L6_L1_FromMinus;
wire MT_Layr_Minus_FM_L5L6_L1_FromMinus_wr_en;
wire [5:0] FM_L5L6_L1_FromMinus_FT_L5L6_number;
wire [9:0] FM_L5L6_L1_FromMinus_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L1_FromMinus_FT_L5L6;
wire FM_L5L6_L1_FromMinus_FT_L5L6_read_en;
FullMatch #(64) FM_L5L6_L1_FromMinus(
.data_in(MT_Layr_Minus_FM_L5L6_L1_FromMinus),
.enable(MT_Layr_Minus_FM_L5L6_L1_FromMinus_wr_en),
.number_out(FM_L5L6_L1_FromMinus_FT_L5L6_number),
.read_add(FM_L5L6_L1_FromMinus_FT_L5L6_read_add),
.data_out(FM_L5L6_L1_FromMinus_FT_L5L6),
.read_en(FM_L5L6_L1_FromMinus_FT_L5L6_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L5L6_L1_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L5L6_L2_FromMinus;
wire MT_Layr_Minus_FM_L5L6_L2_FromMinus_wr_en;
wire [5:0] FM_L5L6_L2_FromMinus_FT_L5L6_number;
wire [9:0] FM_L5L6_L2_FromMinus_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L2_FromMinus_FT_L5L6;
wire FM_L5L6_L2_FromMinus_FT_L5L6_read_en;
FullMatch #(64) FM_L5L6_L2_FromMinus(
.data_in(MT_Layr_Minus_FM_L5L6_L2_FromMinus),
.enable(MT_Layr_Minus_FM_L5L6_L2_FromMinus_wr_en),
.number_out(FM_L5L6_L2_FromMinus_FT_L5L6_number),
.read_add(FM_L5L6_L2_FromMinus_FT_L5L6_read_add),
.data_out(FM_L5L6_L2_FromMinus_FT_L5L6),
.read_en(FM_L5L6_L2_FromMinus_FT_L5L6_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L5L6_L2_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L5L6_L3_FromMinus;
wire MT_Layr_Minus_FM_L5L6_L3_FromMinus_wr_en;
wire [5:0] FM_L5L6_L3_FromMinus_FT_L5L6_number;
wire [9:0] FM_L5L6_L3_FromMinus_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L3_FromMinus_FT_L5L6;
wire FM_L5L6_L3_FromMinus_FT_L5L6_read_en;
FullMatch #(64) FM_L5L6_L3_FromMinus(
.data_in(MT_Layr_Minus_FM_L5L6_L3_FromMinus),
.enable(MT_Layr_Minus_FM_L5L6_L3_FromMinus_wr_en),
.number_out(FM_L5L6_L3_FromMinus_FT_L5L6_number),
.read_add(FM_L5L6_L3_FromMinus_FT_L5L6_read_add),
.data_out(FM_L5L6_L3_FromMinus_FT_L5L6),
.read_en(FM_L5L6_L3_FromMinus_FT_L5L6_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L5L6_L3_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [39:0] MT_Layr_Minus_FM_L5L6_L4_FromMinus;
wire MT_Layr_Minus_FM_L5L6_L4_FromMinus_wr_en;
wire [5:0] FM_L5L6_L4_FromMinus_FT_L5L6_number;
wire [9:0] FM_L5L6_L4_FromMinus_FT_L5L6_read_add;
wire [39:0] FM_L5L6_L4_FromMinus_FT_L5L6;
wire FM_L5L6_L4_FromMinus_FT_L5L6_read_en;
FullMatch #(64) FM_L5L6_L4_FromMinus(
.data_in(MT_Layr_Minus_FM_L5L6_L4_FromMinus),
.enable(MT_Layr_Minus_FM_L5L6_L4_FromMinus_wr_en),
.number_out(FM_L5L6_L4_FromMinus_FT_L5L6_number),
.read_add(FM_L5L6_L4_FromMinus_FT_L5L6_read_add),
.data_out(FM_L5L6_L4_FromMinus_FT_L5L6),
.read_en(FM_L5L6_L4_FromMinus_FT_L5L6_read_en),
.start(MT_Layr_Minus_start),
.done(FM_L5L6_L4_FromMinus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] FT_L1L2_TF_L1L2;
wire FT_L1L2_TF_L1L2_wr_en;
wire [5:0] TF_L1L2_PD_number;
wire [8:0] TF_L1L2_PD_read_add;
wire [125:0] TF_L1L2_PD;
wire [53:0] TF_L1L2_PD_index [`tmux-1:0];
TrackFit  TF_L1L2(
.data_in(FT_L1L2_TF_L1L2),
.enable(FT_L1L2_TF_L1L2_wr_en),
.number_out(TF_L1L2_PD_number),
.read_add(TF_L1L2_PD_read_add),
.data_out(TF_L1L2_PD),
.index_out(TF_L1L2_PD_index),
.start(FT_L1L2_start),
.done(TF_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] FT_L3L4_TF_L3L4;
wire FT_L3L4_TF_L3L4_wr_en;
wire [5:0] TF_L3L4_PD_number;
wire [8:0] TF_L3L4_PD_read_add;
wire [125:0] TF_L3L4_PD;
wire [53:0] TF_L3L4_PD_index [`tmux-1:0];
TrackFit  TF_L3L4(
.data_in(FT_L3L4_TF_L3L4),
.enable(FT_L3L4_TF_L3L4_wr_en),
.number_out(TF_L3L4_PD_number),
.read_add(TF_L3L4_PD_read_add),
.data_out(TF_L3L4_PD),
.index_out(TF_L3L4_PD_index),
.start(FT_L3L4_start),
.done(TF_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] FT_L5L6_TF_L5L6;
wire FT_L5L6_TF_L5L6_wr_en;
wire [5:0] TF_L5L6_PD_number;
wire [8:0] TF_L5L6_PD_read_add;
wire [125:0] TF_L5L6_PD;
wire [53:0] TF_L5L6_PD_index [`tmux-1:0];
TrackFit  TF_L5L6(
.data_in(FT_L5L6_TF_L5L6),
.enable(FT_L5L6_TF_L5L6_wr_en),
.number_out(TF_L5L6_PD_number),
.read_add(TF_L5L6_PD_read_add),
.data_out(TF_L5L6_PD),
.index_out(TF_L5L6_PD_index),
.start(FT_L5L6_start),
.done(TF_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] PD_CT_L1L2;
wire PD_CT_L1L2_wr_en;
//wire CT_L1L2_DataStream;
CleanTrack  CT_L1L2(
.data_in(PD_CT_L1L2),
.enable(PD_CT_L1L2_wr_en),
.data_out(CT_L1L2_DataStream),
.start(PD_start),
.done(CT_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] PD_CT_L3L4;
wire PD_CT_L3L4_wr_en;
//wire CT_L3L4_DataStream;
CleanTrack  CT_L3L4(
.data_in(PD_CT_L3L4),
.enable(PD_CT_L3L4_wr_en),
.data_out(CT_L3L4_DataStream),
.start(PD_start),
.done(CT_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [125:0] PD_CT_L5L6;
wire PD_CT_L5L6_wr_en;
//wire CT_L5L6_DataStream;
CleanTrack  CT_L5L6(
.data_in(PD_CT_L5L6),
.enable(PD_CT_L5L6_wr_en),
.data_out(CT_L5L6_DataStream),
.start(PD_start),
.done(CT_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  LR1_D3(
.stubin(IL1_D3_LR1_D3),
.stubout1(LR1_D3_SL1_L1D3),
.stubout2(LR1_D3_SL1_L2D3),
.stubout3(LR1_D3_SL1_L3D3),
.stubout4(LR1_D3_SL1_L4D3),
.stubout5(LR1_D3_SL1_L5D3),
.stubout6(LR1_D3_SL1_L6D3),
.wr_en1(LR1_D3_SL1_L1D3_wr_en),
.wr_en2(LR1_D3_SL1_L2D3_wr_en),
.wr_en3(LR1_D3_SL1_L3D3_wr_en),
.wr_en4(LR1_D3_SL1_L4D3_wr_en),
.wr_en5(LR1_D3_SL1_L5D3_wr_en),
.wr_en6(LR1_D3_SL1_L6D3_wr_en),
.start(IL1_D3_start),
.done(LR1_D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  LR2_D3(
.stubin(IL2_D3_LR2_D3),
.stubout1(LR2_D3_SL2_L1D3),
.stubout2(LR2_D3_SL2_L2D3),
.stubout3(LR2_D3_SL2_L3D3),
.stubout4(LR2_D3_SL2_L4D3),
.stubout5(LR2_D3_SL2_L5D3),
.stubout6(LR2_D3_SL2_L6D3),
.wr_en1(LR2_D3_SL2_L1D3_wr_en),
.wr_en2(LR2_D3_SL2_L2D3_wr_en),
.wr_en3(LR2_D3_SL2_L3D3_wr_en),
.wr_en4(LR2_D3_SL2_L4D3_wr_en),
.wr_en5(LR2_D3_SL2_L5D3_wr_en),
.wr_en6(LR2_D3_SL2_L6D3_wr_en),
.start(IL2_D3_start),
.done(LR2_D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  LR3_D3(
.stubin(IL3_D3_LR3_D3),
.stubout1(LR3_D3_SL3_L1D3),
.stubout2(LR3_D3_SL3_L2D3),
.stubout3(LR3_D3_SL3_L3D3),
.stubout4(LR3_D3_SL3_L4D3),
.stubout5(LR3_D3_SL3_L5D3),
.stubout6(LR3_D3_SL3_L6D3),
.wr_en1(LR3_D3_SL3_L1D3_wr_en),
.wr_en2(LR3_D3_SL3_L2D3_wr_en),
.wr_en3(LR3_D3_SL3_L3D3_wr_en),
.wr_en4(LR3_D3_SL3_L4D3_wr_en),
.wr_en5(LR3_D3_SL3_L5D3_wr_en),
.wr_en6(LR3_D3_SL3_L6D3_wr_en),
.start(IL3_D3_start),
.done(LR3_D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  LR1_D4(
.stubin(IL1_D4_LR1_D4),
.stubout1(LR1_D4_SL1_L1D4),
.stubout2(LR1_D4_SL1_L2D4),
.stubout3(LR1_D4_SL1_L3D4),
.stubout4(LR1_D4_SL1_L4D4),
.stubout5(LR1_D4_SL1_L5D4),
.stubout6(LR1_D4_SL1_L6D4),
.wr_en1(LR1_D4_SL1_L1D4_wr_en),
.wr_en2(LR1_D4_SL1_L2D4_wr_en),
.wr_en3(LR1_D4_SL1_L3D4_wr_en),
.wr_en4(LR1_D4_SL1_L4D4_wr_en),
.wr_en5(LR1_D4_SL1_L5D4_wr_en),
.wr_en6(LR1_D4_SL1_L6D4_wr_en),
.start(IL1_D4_start),
.done(LR1_D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  LR2_D4(
.stubin(IL2_D4_LR2_D4),
.stubout1(LR2_D4_SL2_L1D4),
.stubout2(LR2_D4_SL2_L2D4),
.stubout3(LR2_D4_SL2_L3D4),
.stubout4(LR2_D4_SL2_L4D4),
.stubout5(LR2_D4_SL2_L5D4),
.stubout6(LR2_D4_SL2_L6D4),
.wr_en1(LR2_D4_SL2_L1D4_wr_en),
.wr_en2(LR2_D4_SL2_L2D4_wr_en),
.wr_en3(LR2_D4_SL2_L3D4_wr_en),
.wr_en4(LR2_D4_SL2_L4D4_wr_en),
.wr_en5(LR2_D4_SL2_L5D4_wr_en),
.wr_en6(LR2_D4_SL2_L6D4_wr_en),
.start(IL2_D4_start),
.done(LR2_D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

LayerRouter  LR3_D4(
.stubin(IL3_D4_LR3_D4),
.stubout1(LR3_D4_SL3_L1D4),
.stubout2(LR3_D4_SL3_L2D4),
.stubout3(LR3_D4_SL3_L3D4),
.stubout4(LR3_D4_SL3_L4D4),
.stubout5(LR3_D4_SL3_L5D4),
.stubout6(LR3_D4_SL3_L6D4),
.wr_en1(LR3_D4_SL3_L1D4_wr_en),
.wr_en2(LR3_D4_SL3_L2D4_wr_en),
.wr_en3(LR3_D4_SL3_L3D4_wr_en),
.wr_en4(LR3_D4_SL3_L4D4_wr_en),
.wr_en5(LR3_D4_SL3_L5D4_wr_en),
.wr_en6(LR3_D4_SL3_L6D4_wr_en),
.start(IL3_D4_start),
.done(LR3_D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b1) VMR_L1D3(
.number_in_stubinLink1(SL1_L1D3_VMR_L1D3_number),
.read_add_stubinLink1(SL1_L1D3_VMR_L1D3_read_add),
.stubinLink1(SL1_L1D3_VMR_L1D3),
.number_in_stubinLink2(SL2_L1D3_VMR_L1D3_number),
.read_add_stubinLink2(SL2_L1D3_VMR_L1D3_read_add),
.stubinLink2(SL2_L1D3_VMR_L1D3),
.number_in_stubinLink3(SL3_L1D3_VMR_L1D3_number),
.read_add_stubinLink3(SL3_L1D3_VMR_L1D3_read_add),
.stubinLink3(SL3_L1D3_VMR_L1D3),
.vmstuboutPHI1X1n1(VMR_L1D3_VMS_L1D3PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L1D3_VMS_L1D3PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L1D3_VMS_L1D3PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L1D3_VMS_L1D3PHI1X1n4),
.vmstuboutPHI1X1n5(VMR_L1D3_VMS_L1D3PHI1X1n5),
.vmstuboutPHI1X1n6(VMR_L1D3_VMS_L1D3PHI1X1n6),
.vmstuboutPHI1X1n7(VMR_L1D3_VMS_L1D3PHI1X1n7),
.vmstuboutPHI1X1n8(VMR_L1D3_VMS_L1D3PHI1X1n8),
.vmstuboutPHI2X1n1(VMR_L1D3_VMS_L1D3PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L1D3_VMS_L1D3PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L1D3_VMS_L1D3PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L1D3_VMS_L1D3PHI2X1n4),
.vmstuboutPHI2X1n5(VMR_L1D3_VMS_L1D3PHI2X1n5),
.vmstuboutPHI2X1n6(VMR_L1D3_VMS_L1D3PHI2X1n6),
.vmstuboutPHI2X1n7(VMR_L1D3_VMS_L1D3PHI2X1n7),
.vmstuboutPHI2X1n8(VMR_L1D3_VMS_L1D3PHI2X1n8),
.vmstuboutPHI3X1n1(VMR_L1D3_VMS_L1D3PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L1D3_VMS_L1D3PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L1D3_VMS_L1D3PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L1D3_VMS_L1D3PHI3X1n4),
.vmstuboutPHI3X1n5(VMR_L1D3_VMS_L1D3PHI3X1n5),
.vmstuboutPHI3X1n6(VMR_L1D3_VMS_L1D3PHI3X1n6),
.vmstuboutPHI3X1n7(VMR_L1D3_VMS_L1D3PHI3X1n7),
.vmstuboutPHI3X1n8(VMR_L1D3_VMS_L1D3PHI3X1n8),
.vmstuboutPHI1X2n1(VMR_L1D3_VMS_L1D3PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L1D3_VMS_L1D3PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L1D3_VMS_L1D3PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L1D3_VMS_L1D3PHI1X2n4),
.vmstuboutPHI1X2n5(VMR_L1D3_VMS_L1D3PHI1X2n5),
.vmstuboutPHI1X2n6(VMR_L1D3_VMS_L1D3PHI1X2n6),
.vmstuboutPHI1X2n7(VMR_L1D3_VMS_L1D3PHI1X2n7),
.vmstuboutPHI1X2n8(VMR_L1D3_VMS_L1D3PHI1X2n8),
.vmstuboutPHI2X2n1(VMR_L1D3_VMS_L1D3PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L1D3_VMS_L1D3PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L1D3_VMS_L1D3PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L1D3_VMS_L1D3PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L1D3_VMS_L1D3PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L1D3_VMS_L1D3PHI2X2n6),
.vmstuboutPHI2X2n7(VMR_L1D3_VMS_L1D3PHI2X2n7),
.vmstuboutPHI2X2n8(VMR_L1D3_VMS_L1D3PHI2X2n8),
.vmstuboutPHI3X2n1(VMR_L1D3_VMS_L1D3PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L1D3_VMS_L1D3PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L1D3_VMS_L1D3PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L1D3_VMS_L1D3PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L1D3_VMS_L1D3PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L1D3_VMS_L1D3PHI3X2n6),
.vmstuboutPHI3X2n7(VMR_L1D3_VMS_L1D3PHI3X2n7),
.vmstuboutPHI3X2n8(VMR_L1D3_VMS_L1D3PHI3X2n8),
.allstuboutn1(VMR_L1D3_AS_L1D3n1),
.allstuboutn2(VMR_L1D3_AS_L1D3n2),
.allstuboutn3(VMR_L1D3_AS_L1D3n3),
.allstuboutn4(VMR_L1D3_AS_L1D3n4),
.vmstuboutPHI1X1n1_wr_en(VMR_L1D3_VMS_L1D3PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L1D3_VMS_L1D3PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L1D3_VMS_L1D3PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L1D3_VMS_L1D3PHI1X1n4_wr_en),
.vmstuboutPHI1X1n5_wr_en(VMR_L1D3_VMS_L1D3PHI1X1n5_wr_en),
.vmstuboutPHI1X1n6_wr_en(VMR_L1D3_VMS_L1D3PHI1X1n6_wr_en),
.vmstuboutPHI1X1n7_wr_en(VMR_L1D3_VMS_L1D3PHI1X1n7_wr_en),
.vmstuboutPHI1X1n8_wr_en(VMR_L1D3_VMS_L1D3PHI1X1n8_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L1D3_VMS_L1D3PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L1D3_VMS_L1D3PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L1D3_VMS_L1D3PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L1D3_VMS_L1D3PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMR_L1D3_VMS_L1D3PHI2X1n5_wr_en),
.vmstuboutPHI2X1n6_wr_en(VMR_L1D3_VMS_L1D3PHI2X1n6_wr_en),
.vmstuboutPHI2X1n7_wr_en(VMR_L1D3_VMS_L1D3PHI2X1n7_wr_en),
.vmstuboutPHI2X1n8_wr_en(VMR_L1D3_VMS_L1D3PHI2X1n8_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L1D3_VMS_L1D3PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L1D3_VMS_L1D3PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L1D3_VMS_L1D3PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L1D3_VMS_L1D3PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMR_L1D3_VMS_L1D3PHI3X1n5_wr_en),
.vmstuboutPHI3X1n6_wr_en(VMR_L1D3_VMS_L1D3PHI3X1n6_wr_en),
.vmstuboutPHI3X1n7_wr_en(VMR_L1D3_VMS_L1D3PHI3X1n7_wr_en),
.vmstuboutPHI3X1n8_wr_en(VMR_L1D3_VMS_L1D3PHI3X1n8_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L1D3_VMS_L1D3PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L1D3_VMS_L1D3PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L1D3_VMS_L1D3PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L1D3_VMS_L1D3PHI1X2n4_wr_en),
.vmstuboutPHI1X2n5_wr_en(VMR_L1D3_VMS_L1D3PHI1X2n5_wr_en),
.vmstuboutPHI1X2n6_wr_en(VMR_L1D3_VMS_L1D3PHI1X2n6_wr_en),
.vmstuboutPHI1X2n7_wr_en(VMR_L1D3_VMS_L1D3PHI1X2n7_wr_en),
.vmstuboutPHI1X2n8_wr_en(VMR_L1D3_VMS_L1D3PHI1X2n8_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L1D3_VMS_L1D3PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L1D3_VMS_L1D3PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L1D3_VMS_L1D3PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L1D3_VMS_L1D3PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L1D3_VMS_L1D3PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L1D3_VMS_L1D3PHI2X2n6_wr_en),
.vmstuboutPHI2X2n7_wr_en(VMR_L1D3_VMS_L1D3PHI2X2n7_wr_en),
.vmstuboutPHI2X2n8_wr_en(VMR_L1D3_VMS_L1D3PHI2X2n8_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L1D3_VMS_L1D3PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L1D3_VMS_L1D3PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L1D3_VMS_L1D3PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L1D3_VMS_L1D3PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L1D3_VMS_L1D3PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L1D3_VMS_L1D3PHI3X2n6_wr_en),
.vmstuboutPHI3X2n7_wr_en(VMR_L1D3_VMS_L1D3PHI3X2n7_wr_en),
.vmstuboutPHI3X2n8_wr_en(VMR_L1D3_VMS_L1D3PHI3X2n8_wr_en),
.valid_data1(VMR_L1D3_AS_L1D3n1_wr_en),
.valid_data2(VMR_L1D3_AS_L1D3n2_wr_en),
.valid_data3(VMR_L1D3_AS_L1D3n3_wr_en),
.valid_data4(VMR_L1D3_AS_L1D3n4_wr_en),
.start(SL1_L1D3_start),
.done(VMR_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b1) VMR_L1D4(
.number_in_stubinLink1(SL1_L1D4_VMR_L1D4_number),
.read_add_stubinLink1(SL1_L1D4_VMR_L1D4_read_add),
.stubinLink1(SL1_L1D4_VMR_L1D4),
.number_in_stubinLink2(SL2_L1D4_VMR_L1D4_number),
.read_add_stubinLink2(SL2_L1D4_VMR_L1D4_read_add),
.stubinLink2(SL2_L1D4_VMR_L1D4),
.number_in_stubinLink3(SL3_L1D4_VMR_L1D4_number),
.read_add_stubinLink3(SL3_L1D4_VMR_L1D4_read_add),
.stubinLink3(SL3_L1D4_VMR_L1D4),
.vmstuboutPHI1X1n1(VMR_L1D4_VMS_L1D4PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L1D4_VMS_L1D4PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L1D4_VMS_L1D4PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L1D4_VMS_L1D4PHI1X1n4),
.vmstuboutPHI2X1n1(VMR_L1D4_VMS_L1D4PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L1D4_VMS_L1D4PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L1D4_VMS_L1D4PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L1D4_VMS_L1D4PHI2X1n4),
.vmstuboutPHI3X1n1(VMR_L1D4_VMS_L1D4PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L1D4_VMS_L1D4PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L1D4_VMS_L1D4PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L1D4_VMS_L1D4PHI3X1n4),
.allstuboutn1(VMR_L1D4_AS_L1D4n1),
.allstuboutn2(VMR_L1D4_AS_L1D4n2),
.allstuboutn3(VMR_L1D4_AS_L1D4n3),
.vmstuboutPHI1X2n1(VMR_L1D4_VMS_L1D4PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L1D4_VMS_L1D4PHI1X2n2),
.vmstuboutPHI2X2n1(VMR_L1D4_VMS_L1D4PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L1D4_VMS_L1D4PHI2X2n2),
.vmstuboutPHI3X2n1(VMR_L1D4_VMS_L1D4PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L1D4_VMS_L1D4PHI3X2n2),
.vmstuboutPHI1X1n1_wr_en(VMR_L1D4_VMS_L1D4PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L1D4_VMS_L1D4PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L1D4_VMS_L1D4PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L1D4_VMS_L1D4PHI1X1n4_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L1D4_VMS_L1D4PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L1D4_VMS_L1D4PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L1D4_VMS_L1D4PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L1D4_VMS_L1D4PHI2X1n4_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L1D4_VMS_L1D4PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L1D4_VMS_L1D4PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L1D4_VMS_L1D4PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L1D4_VMS_L1D4PHI3X1n4_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L1D4_VMS_L1D4PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L1D4_VMS_L1D4PHI1X2n2_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L1D4_VMS_L1D4PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L1D4_VMS_L1D4PHI2X2n2_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L1D4_VMS_L1D4PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L1D4_VMS_L1D4PHI3X2n2_wr_en),
.valid_data1(VMR_L1D4_AS_L1D4n1_wr_en),
.valid_data2(VMR_L1D4_AS_L1D4n2_wr_en),
.valid_data3(VMR_L1D4_AS_L1D4n3_wr_en),
.start(SL1_L1D4_start),
.done(VMR_L1D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b0) VMR_L2D3(
.number_in_stubinLink1(SL1_L2D3_VMR_L2D3_number),
.read_add_stubinLink1(SL1_L2D3_VMR_L2D3_read_add),
.stubinLink1(SL1_L2D3_VMR_L2D3),
.number_in_stubinLink2(SL2_L2D3_VMR_L2D3_number),
.read_add_stubinLink2(SL2_L2D3_VMR_L2D3_read_add),
.stubinLink2(SL2_L2D3_VMR_L2D3),
.number_in_stubinLink3(SL3_L2D3_VMR_L2D3_number),
.read_add_stubinLink3(SL3_L2D3_VMR_L2D3_read_add),
.stubinLink3(SL3_L2D3_VMR_L2D3),
.vmstuboutPHI1X1n1(VMR_L2D3_VMS_L2D3PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L2D3_VMS_L2D3PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L2D3_VMS_L2D3PHI1X1n3),
.vmstuboutPHI2X1n1(VMR_L2D3_VMS_L2D3PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L2D3_VMS_L2D3PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L2D3_VMS_L2D3PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L2D3_VMS_L2D3PHI2X1n4),
.vmstuboutPHI3X1n1(VMR_L2D3_VMS_L2D3PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L2D3_VMS_L2D3PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L2D3_VMS_L2D3PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L2D3_VMS_L2D3PHI3X1n4),
.vmstuboutPHI4X1n1(VMR_L2D3_VMS_L2D3PHI4X1n1),
.vmstuboutPHI4X1n2(VMR_L2D3_VMS_L2D3PHI4X1n2),
.vmstuboutPHI4X1n3(VMR_L2D3_VMS_L2D3PHI4X1n3),
.vmstuboutPHI1X2n1(VMR_L2D3_VMS_L2D3PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L2D3_VMS_L2D3PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L2D3_VMS_L2D3PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L2D3_VMS_L2D3PHI1X2n4),
.vmstuboutPHI2X2n1(VMR_L2D3_VMS_L2D3PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L2D3_VMS_L2D3PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L2D3_VMS_L2D3PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L2D3_VMS_L2D3PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L2D3_VMS_L2D3PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L2D3_VMS_L2D3PHI2X2n6),
.vmstuboutPHI3X2n1(VMR_L2D3_VMS_L2D3PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L2D3_VMS_L2D3PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L2D3_VMS_L2D3PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L2D3_VMS_L2D3PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L2D3_VMS_L2D3PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L2D3_VMS_L2D3PHI3X2n6),
.vmstuboutPHI4X2n1(VMR_L2D3_VMS_L2D3PHI4X2n1),
.vmstuboutPHI4X2n2(VMR_L2D3_VMS_L2D3PHI4X2n2),
.vmstuboutPHI4X2n3(VMR_L2D3_VMS_L2D3PHI4X2n3),
.vmstuboutPHI4X2n4(VMR_L2D3_VMS_L2D3PHI4X2n4),
.allstuboutn1(VMR_L2D3_AS_L2D3n1),
.allstuboutn2(VMR_L2D3_AS_L2D3n2),
.allstuboutn3(VMR_L2D3_AS_L2D3n3),
.vmstuboutPHI1X1n1_wr_en(VMR_L2D3_VMS_L2D3PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L2D3_VMS_L2D3PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L2D3_VMS_L2D3PHI1X1n3_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L2D3_VMS_L2D3PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L2D3_VMS_L2D3PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L2D3_VMS_L2D3PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L2D3_VMS_L2D3PHI2X1n4_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L2D3_VMS_L2D3PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L2D3_VMS_L2D3PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L2D3_VMS_L2D3PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L2D3_VMS_L2D3PHI3X1n4_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMR_L2D3_VMS_L2D3PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMR_L2D3_VMS_L2D3PHI4X1n2_wr_en),
.vmstuboutPHI4X1n3_wr_en(VMR_L2D3_VMS_L2D3PHI4X1n3_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L2D3_VMS_L2D3PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L2D3_VMS_L2D3PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L2D3_VMS_L2D3PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L2D3_VMS_L2D3PHI1X2n4_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L2D3_VMS_L2D3PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L2D3_VMS_L2D3PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L2D3_VMS_L2D3PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L2D3_VMS_L2D3PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L2D3_VMS_L2D3PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L2D3_VMS_L2D3PHI2X2n6_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L2D3_VMS_L2D3PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L2D3_VMS_L2D3PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L2D3_VMS_L2D3PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L2D3_VMS_L2D3PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L2D3_VMS_L2D3PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L2D3_VMS_L2D3PHI3X2n6_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMR_L2D3_VMS_L2D3PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMR_L2D3_VMS_L2D3PHI4X2n2_wr_en),
.vmstuboutPHI4X2n3_wr_en(VMR_L2D3_VMS_L2D3PHI4X2n3_wr_en),
.vmstuboutPHI4X2n4_wr_en(VMR_L2D3_VMS_L2D3PHI4X2n4_wr_en),
.valid_data1(VMR_L2D3_AS_L2D3n1_wr_en),
.valid_data2(VMR_L2D3_AS_L2D3n2_wr_en),
.valid_data3(VMR_L2D3_AS_L2D3n3_wr_en),
.start(SL1_L2D3_start),
.done(VMR_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b0) VMR_L2D4(
.number_in_stubinLink1(SL1_L2D4_VMR_L2D4_number),
.read_add_stubinLink1(SL1_L2D4_VMR_L2D4_read_add),
.stubinLink1(SL1_L2D4_VMR_L2D4),
.number_in_stubinLink2(SL2_L2D4_VMR_L2D4_number),
.read_add_stubinLink2(SL2_L2D4_VMR_L2D4_read_add),
.stubinLink2(SL2_L2D4_VMR_L2D4),
.number_in_stubinLink3(SL3_L2D4_VMR_L2D4_number),
.read_add_stubinLink3(SL3_L2D4_VMR_L2D4_read_add),
.stubinLink3(SL3_L2D4_VMR_L2D4),
.vmstuboutPHI1X1n1(VMR_L2D4_VMS_L2D4PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L2D4_VMS_L2D4PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L2D4_VMS_L2D4PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L2D4_VMS_L2D4PHI1X1n4),
.vmstuboutPHI2X1n1(VMR_L2D4_VMS_L2D4PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L2D4_VMS_L2D4PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L2D4_VMS_L2D4PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L2D4_VMS_L2D4PHI2X1n4),
.vmstuboutPHI2X1n5(VMR_L2D4_VMS_L2D4PHI2X1n5),
.vmstuboutPHI2X1n6(VMR_L2D4_VMS_L2D4PHI2X1n6),
.vmstuboutPHI3X1n1(VMR_L2D4_VMS_L2D4PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L2D4_VMS_L2D4PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L2D4_VMS_L2D4PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L2D4_VMS_L2D4PHI3X1n4),
.vmstuboutPHI3X1n5(VMR_L2D4_VMS_L2D4PHI3X1n5),
.vmstuboutPHI3X1n6(VMR_L2D4_VMS_L2D4PHI3X1n6),
.vmstuboutPHI4X1n1(VMR_L2D4_VMS_L2D4PHI4X1n1),
.vmstuboutPHI4X1n2(VMR_L2D4_VMS_L2D4PHI4X1n2),
.vmstuboutPHI4X1n3(VMR_L2D4_VMS_L2D4PHI4X1n3),
.vmstuboutPHI4X1n4(VMR_L2D4_VMS_L2D4PHI4X1n4),
.vmstuboutPHI1X2n1(VMR_L2D4_VMS_L2D4PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L2D4_VMS_L2D4PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L2D4_VMS_L2D4PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L2D4_VMS_L2D4PHI1X2n4),
.vmstuboutPHI2X2n1(VMR_L2D4_VMS_L2D4PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L2D4_VMS_L2D4PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L2D4_VMS_L2D4PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L2D4_VMS_L2D4PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L2D4_VMS_L2D4PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L2D4_VMS_L2D4PHI2X2n6),
.vmstuboutPHI3X2n1(VMR_L2D4_VMS_L2D4PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L2D4_VMS_L2D4PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L2D4_VMS_L2D4PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L2D4_VMS_L2D4PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L2D4_VMS_L2D4PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L2D4_VMS_L2D4PHI3X2n6),
.vmstuboutPHI4X2n1(VMR_L2D4_VMS_L2D4PHI4X2n1),
.vmstuboutPHI4X2n2(VMR_L2D4_VMS_L2D4PHI4X2n2),
.vmstuboutPHI4X2n3(VMR_L2D4_VMS_L2D4PHI4X2n3),
.vmstuboutPHI4X2n4(VMR_L2D4_VMS_L2D4PHI4X2n4),
.allstuboutn1(VMR_L2D4_AS_L2D4n1),
.allstuboutn2(VMR_L2D4_AS_L2D4n2),
.allstuboutn3(VMR_L2D4_AS_L2D4n3),
.allstuboutn4(VMR_L2D4_AS_L2D4n4),
.vmstuboutPHI1X1n1_wr_en(VMR_L2D4_VMS_L2D4PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L2D4_VMS_L2D4PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L2D4_VMS_L2D4PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L2D4_VMS_L2D4PHI1X1n4_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L2D4_VMS_L2D4PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L2D4_VMS_L2D4PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L2D4_VMS_L2D4PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L2D4_VMS_L2D4PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMR_L2D4_VMS_L2D4PHI2X1n5_wr_en),
.vmstuboutPHI2X1n6_wr_en(VMR_L2D4_VMS_L2D4PHI2X1n6_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L2D4_VMS_L2D4PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L2D4_VMS_L2D4PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L2D4_VMS_L2D4PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L2D4_VMS_L2D4PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMR_L2D4_VMS_L2D4PHI3X1n5_wr_en),
.vmstuboutPHI3X1n6_wr_en(VMR_L2D4_VMS_L2D4PHI3X1n6_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMR_L2D4_VMS_L2D4PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMR_L2D4_VMS_L2D4PHI4X1n2_wr_en),
.vmstuboutPHI4X1n3_wr_en(VMR_L2D4_VMS_L2D4PHI4X1n3_wr_en),
.vmstuboutPHI4X1n4_wr_en(VMR_L2D4_VMS_L2D4PHI4X1n4_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L2D4_VMS_L2D4PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L2D4_VMS_L2D4PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L2D4_VMS_L2D4PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L2D4_VMS_L2D4PHI1X2n4_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L2D4_VMS_L2D4PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L2D4_VMS_L2D4PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L2D4_VMS_L2D4PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L2D4_VMS_L2D4PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L2D4_VMS_L2D4PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L2D4_VMS_L2D4PHI2X2n6_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L2D4_VMS_L2D4PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L2D4_VMS_L2D4PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L2D4_VMS_L2D4PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L2D4_VMS_L2D4PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L2D4_VMS_L2D4PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L2D4_VMS_L2D4PHI3X2n6_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMR_L2D4_VMS_L2D4PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMR_L2D4_VMS_L2D4PHI4X2n2_wr_en),
.vmstuboutPHI4X2n3_wr_en(VMR_L2D4_VMS_L2D4PHI4X2n3_wr_en),
.vmstuboutPHI4X2n4_wr_en(VMR_L2D4_VMS_L2D4PHI4X2n4_wr_en),
.valid_data1(VMR_L2D4_AS_L2D4n1_wr_en),
.valid_data2(VMR_L2D4_AS_L2D4n2_wr_en),
.valid_data3(VMR_L2D4_AS_L2D4n3_wr_en),
.valid_data4(VMR_L2D4_AS_L2D4n4_wr_en),
.start(SL1_L2D4_start),
.done(VMR_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b1) VMR_L3D3(
.number_in_stubinLink1(SL1_L3D3_VMR_L3D3_number),
.read_add_stubinLink1(SL1_L3D3_VMR_L3D3_read_add),
.stubinLink1(SL1_L3D3_VMR_L3D3),
.number_in_stubinLink2(SL2_L3D3_VMR_L3D3_number),
.read_add_stubinLink2(SL2_L3D3_VMR_L3D3_read_add),
.stubinLink2(SL2_L3D3_VMR_L3D3),
.number_in_stubinLink3(SL3_L3D3_VMR_L3D3_number),
.read_add_stubinLink3(SL3_L3D3_VMR_L3D3_read_add),
.stubinLink3(SL3_L3D3_VMR_L3D3),
.vmstuboutPHI1X1n1(VMR_L3D3_VMS_L3D3PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L3D3_VMS_L3D3PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L3D3_VMS_L3D3PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L3D3_VMS_L3D3PHI1X1n4),
.vmstuboutPHI1X1n5(VMR_L3D3_VMS_L3D3PHI1X1n5),
.vmstuboutPHI1X1n6(VMR_L3D3_VMS_L3D3PHI1X1n6),
.vmstuboutPHI2X1n1(VMR_L3D3_VMS_L3D3PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L3D3_VMS_L3D3PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L3D3_VMS_L3D3PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L3D3_VMS_L3D3PHI2X1n4),
.vmstuboutPHI2X1n5(VMR_L3D3_VMS_L3D3PHI2X1n5),
.vmstuboutPHI2X1n6(VMR_L3D3_VMS_L3D3PHI2X1n6),
.vmstuboutPHI3X1n1(VMR_L3D3_VMS_L3D3PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L3D3_VMS_L3D3PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L3D3_VMS_L3D3PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L3D3_VMS_L3D3PHI3X1n4),
.vmstuboutPHI3X1n5(VMR_L3D3_VMS_L3D3PHI3X1n5),
.vmstuboutPHI3X1n6(VMR_L3D3_VMS_L3D3PHI3X1n6),
.vmstuboutPHI1X2n1(VMR_L3D3_VMS_L3D3PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L3D3_VMS_L3D3PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L3D3_VMS_L3D3PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L3D3_VMS_L3D3PHI1X2n4),
.vmstuboutPHI1X2n5(VMR_L3D3_VMS_L3D3PHI1X2n5),
.vmstuboutPHI1X2n6(VMR_L3D3_VMS_L3D3PHI1X2n6),
.vmstuboutPHI2X2n1(VMR_L3D3_VMS_L3D3PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L3D3_VMS_L3D3PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L3D3_VMS_L3D3PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L3D3_VMS_L3D3PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L3D3_VMS_L3D3PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L3D3_VMS_L3D3PHI2X2n6),
.vmstuboutPHI3X2n1(VMR_L3D3_VMS_L3D3PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L3D3_VMS_L3D3PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L3D3_VMS_L3D3PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L3D3_VMS_L3D3PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L3D3_VMS_L3D3PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L3D3_VMS_L3D3PHI3X2n6),
.allstuboutn1(VMR_L3D3_AS_L3D3n1),
.allstuboutn2(VMR_L3D3_AS_L3D3n2),
.allstuboutn3(VMR_L3D3_AS_L3D3n3),
.allstuboutn4(VMR_L3D3_AS_L3D3n4),
.vmstuboutPHI1X1n1_wr_en(VMR_L3D3_VMS_L3D3PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L3D3_VMS_L3D3PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L3D3_VMS_L3D3PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L3D3_VMS_L3D3PHI1X1n4_wr_en),
.vmstuboutPHI1X1n5_wr_en(VMR_L3D3_VMS_L3D3PHI1X1n5_wr_en),
.vmstuboutPHI1X1n6_wr_en(VMR_L3D3_VMS_L3D3PHI1X1n6_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L3D3_VMS_L3D3PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L3D3_VMS_L3D3PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L3D3_VMS_L3D3PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L3D3_VMS_L3D3PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMR_L3D3_VMS_L3D3PHI2X1n5_wr_en),
.vmstuboutPHI2X1n6_wr_en(VMR_L3D3_VMS_L3D3PHI2X1n6_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L3D3_VMS_L3D3PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L3D3_VMS_L3D3PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L3D3_VMS_L3D3PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L3D3_VMS_L3D3PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMR_L3D3_VMS_L3D3PHI3X1n5_wr_en),
.vmstuboutPHI3X1n6_wr_en(VMR_L3D3_VMS_L3D3PHI3X1n6_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L3D3_VMS_L3D3PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L3D3_VMS_L3D3PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L3D3_VMS_L3D3PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L3D3_VMS_L3D3PHI1X2n4_wr_en),
.vmstuboutPHI1X2n5_wr_en(VMR_L3D3_VMS_L3D3PHI1X2n5_wr_en),
.vmstuboutPHI1X2n6_wr_en(VMR_L3D3_VMS_L3D3PHI1X2n6_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L3D3_VMS_L3D3PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L3D3_VMS_L3D3PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L3D3_VMS_L3D3PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L3D3_VMS_L3D3PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L3D3_VMS_L3D3PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L3D3_VMS_L3D3PHI2X2n6_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L3D3_VMS_L3D3PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L3D3_VMS_L3D3PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L3D3_VMS_L3D3PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L3D3_VMS_L3D3PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L3D3_VMS_L3D3PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L3D3_VMS_L3D3PHI3X2n6_wr_en),
.valid_data1(VMR_L3D3_AS_L3D3n1_wr_en),
.valid_data2(VMR_L3D3_AS_L3D3n2_wr_en),
.valid_data3(VMR_L3D3_AS_L3D3n3_wr_en),
.valid_data4(VMR_L3D3_AS_L3D3n4_wr_en),
.start(SL1_L3D3_start),
.done(VMR_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b1,1'b1) VMR_L3D4(
.number_in_stubinLink1(SL1_L3D4_VMR_L3D4_number),
.read_add_stubinLink1(SL1_L3D4_VMR_L3D4_read_add),
.stubinLink1(SL1_L3D4_VMR_L3D4),
.number_in_stubinLink2(SL2_L3D4_VMR_L3D4_number),
.read_add_stubinLink2(SL2_L3D4_VMR_L3D4_read_add),
.stubinLink2(SL2_L3D4_VMR_L3D4),
.number_in_stubinLink3(SL3_L3D4_VMR_L3D4_number),
.read_add_stubinLink3(SL3_L3D4_VMR_L3D4_read_add),
.stubinLink3(SL3_L3D4_VMR_L3D4),
.vmstuboutPHI1X1n1(VMR_L3D4_VMS_L3D4PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L3D4_VMS_L3D4PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L3D4_VMS_L3D4PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L3D4_VMS_L3D4PHI1X1n4),
.vmstuboutPHI1X1n5(VMR_L3D4_VMS_L3D4PHI1X1n5),
.vmstuboutPHI1X1n6(VMR_L3D4_VMS_L3D4PHI1X1n6),
.vmstuboutPHI2X1n1(VMR_L3D4_VMS_L3D4PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L3D4_VMS_L3D4PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L3D4_VMS_L3D4PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L3D4_VMS_L3D4PHI2X1n4),
.vmstuboutPHI2X1n5(VMR_L3D4_VMS_L3D4PHI2X1n5),
.vmstuboutPHI2X1n6(VMR_L3D4_VMS_L3D4PHI2X1n6),
.vmstuboutPHI3X1n1(VMR_L3D4_VMS_L3D4PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L3D4_VMS_L3D4PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L3D4_VMS_L3D4PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L3D4_VMS_L3D4PHI3X1n4),
.vmstuboutPHI3X1n5(VMR_L3D4_VMS_L3D4PHI3X1n5),
.vmstuboutPHI3X1n6(VMR_L3D4_VMS_L3D4PHI3X1n6),
.vmstuboutPHI1X2n1(VMR_L3D4_VMS_L3D4PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L3D4_VMS_L3D4PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L3D4_VMS_L3D4PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L3D4_VMS_L3D4PHI1X2n4),
.vmstuboutPHI2X2n1(VMR_L3D4_VMS_L3D4PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L3D4_VMS_L3D4PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L3D4_VMS_L3D4PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L3D4_VMS_L3D4PHI2X2n4),
.vmstuboutPHI3X2n1(VMR_L3D4_VMS_L3D4PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L3D4_VMS_L3D4PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L3D4_VMS_L3D4PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L3D4_VMS_L3D4PHI3X2n4),
.allstuboutn1(VMR_L3D4_AS_L3D4n1),
.allstuboutn2(VMR_L3D4_AS_L3D4n2),
.allstuboutn3(VMR_L3D4_AS_L3D4n3),
.vmstuboutPHI1X1n1_wr_en(VMR_L3D4_VMS_L3D4PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L3D4_VMS_L3D4PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L3D4_VMS_L3D4PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L3D4_VMS_L3D4PHI1X1n4_wr_en),
.vmstuboutPHI1X1n5_wr_en(VMR_L3D4_VMS_L3D4PHI1X1n5_wr_en),
.vmstuboutPHI1X1n6_wr_en(VMR_L3D4_VMS_L3D4PHI1X1n6_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L3D4_VMS_L3D4PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L3D4_VMS_L3D4PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L3D4_VMS_L3D4PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L3D4_VMS_L3D4PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMR_L3D4_VMS_L3D4PHI2X1n5_wr_en),
.vmstuboutPHI2X1n6_wr_en(VMR_L3D4_VMS_L3D4PHI2X1n6_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L3D4_VMS_L3D4PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L3D4_VMS_L3D4PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L3D4_VMS_L3D4PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L3D4_VMS_L3D4PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMR_L3D4_VMS_L3D4PHI3X1n5_wr_en),
.vmstuboutPHI3X1n6_wr_en(VMR_L3D4_VMS_L3D4PHI3X1n6_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L3D4_VMS_L3D4PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L3D4_VMS_L3D4PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L3D4_VMS_L3D4PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L3D4_VMS_L3D4PHI1X2n4_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L3D4_VMS_L3D4PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L3D4_VMS_L3D4PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L3D4_VMS_L3D4PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L3D4_VMS_L3D4PHI2X2n4_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L3D4_VMS_L3D4PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L3D4_VMS_L3D4PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L3D4_VMS_L3D4PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L3D4_VMS_L3D4PHI3X2n4_wr_en),
.valid_data1(VMR_L3D4_AS_L3D4n1_wr_en),
.valid_data2(VMR_L3D4_AS_L3D4n2_wr_en),
.valid_data3(VMR_L3D4_AS_L3D4n3_wr_en),
.start(SL1_L3D4_start),
.done(VMR_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b0,1'b0) VMR_L4D3(
.number_in_stubinLink1(SL1_L4D3_VMR_L4D3_number),
.read_add_stubinLink1(SL1_L4D3_VMR_L4D3_read_add),
.stubinLink1(SL1_L4D3_VMR_L4D3),
.number_in_stubinLink2(SL2_L4D3_VMR_L4D3_number),
.read_add_stubinLink2(SL2_L4D3_VMR_L4D3_read_add),
.stubinLink2(SL2_L4D3_VMR_L4D3),
.number_in_stubinLink3(SL3_L4D3_VMR_L4D3_number),
.read_add_stubinLink3(SL3_L4D3_VMR_L4D3_read_add),
.stubinLink3(SL3_L4D3_VMR_L4D3),
.vmstuboutPHI1X1n1(VMR_L4D3_VMS_L4D3PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L4D3_VMS_L4D3PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L4D3_VMS_L4D3PHI1X1n3),
.vmstuboutPHI2X1n1(VMR_L4D3_VMS_L4D3PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L4D3_VMS_L4D3PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L4D3_VMS_L4D3PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L4D3_VMS_L4D3PHI2X1n4),
.vmstuboutPHI3X1n1(VMR_L4D3_VMS_L4D3PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L4D3_VMS_L4D3PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L4D3_VMS_L4D3PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L4D3_VMS_L4D3PHI3X1n4),
.vmstuboutPHI4X1n1(VMR_L4D3_VMS_L4D3PHI4X1n1),
.vmstuboutPHI4X1n2(VMR_L4D3_VMS_L4D3PHI4X1n2),
.vmstuboutPHI4X1n3(VMR_L4D3_VMS_L4D3PHI4X1n3),
.vmstuboutPHI1X2n1(VMR_L4D3_VMS_L4D3PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L4D3_VMS_L4D3PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L4D3_VMS_L4D3PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L4D3_VMS_L4D3PHI1X2n4),
.vmstuboutPHI2X2n1(VMR_L4D3_VMS_L4D3PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L4D3_VMS_L4D3PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L4D3_VMS_L4D3PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L4D3_VMS_L4D3PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L4D3_VMS_L4D3PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L4D3_VMS_L4D3PHI2X2n6),
.vmstuboutPHI3X2n1(VMR_L4D3_VMS_L4D3PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L4D3_VMS_L4D3PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L4D3_VMS_L4D3PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L4D3_VMS_L4D3PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L4D3_VMS_L4D3PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L4D3_VMS_L4D3PHI3X2n6),
.vmstuboutPHI4X2n1(VMR_L4D3_VMS_L4D3PHI4X2n1),
.vmstuboutPHI4X2n2(VMR_L4D3_VMS_L4D3PHI4X2n2),
.vmstuboutPHI4X2n3(VMR_L4D3_VMS_L4D3PHI4X2n3),
.vmstuboutPHI4X2n4(VMR_L4D3_VMS_L4D3PHI4X2n4),
.allstuboutn1(VMR_L4D3_AS_L4D3n1),
.allstuboutn2(VMR_L4D3_AS_L4D3n2),
.allstuboutn3(VMR_L4D3_AS_L4D3n3),
.vmstuboutPHI1X1n1_wr_en(VMR_L4D3_VMS_L4D3PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L4D3_VMS_L4D3PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L4D3_VMS_L4D3PHI1X1n3_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L4D3_VMS_L4D3PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L4D3_VMS_L4D3PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L4D3_VMS_L4D3PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L4D3_VMS_L4D3PHI2X1n4_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L4D3_VMS_L4D3PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L4D3_VMS_L4D3PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L4D3_VMS_L4D3PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L4D3_VMS_L4D3PHI3X1n4_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMR_L4D3_VMS_L4D3PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMR_L4D3_VMS_L4D3PHI4X1n2_wr_en),
.vmstuboutPHI4X1n3_wr_en(VMR_L4D3_VMS_L4D3PHI4X1n3_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L4D3_VMS_L4D3PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L4D3_VMS_L4D3PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L4D3_VMS_L4D3PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L4D3_VMS_L4D3PHI1X2n4_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L4D3_VMS_L4D3PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L4D3_VMS_L4D3PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L4D3_VMS_L4D3PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L4D3_VMS_L4D3PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L4D3_VMS_L4D3PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L4D3_VMS_L4D3PHI2X2n6_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L4D3_VMS_L4D3PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L4D3_VMS_L4D3PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L4D3_VMS_L4D3PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L4D3_VMS_L4D3PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L4D3_VMS_L4D3PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L4D3_VMS_L4D3PHI3X2n6_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMR_L4D3_VMS_L4D3PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMR_L4D3_VMS_L4D3PHI4X2n2_wr_en),
.vmstuboutPHI4X2n3_wr_en(VMR_L4D3_VMS_L4D3PHI4X2n3_wr_en),
.vmstuboutPHI4X2n4_wr_en(VMR_L4D3_VMS_L4D3PHI4X2n4_wr_en),
.valid_data1(VMR_L4D3_AS_L4D3n1_wr_en),
.valid_data2(VMR_L4D3_AS_L4D3n2_wr_en),
.valid_data3(VMR_L4D3_AS_L4D3n3_wr_en),
.start(SL1_L4D3_start),
.done(VMR_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b0,1'b0) VMR_L4D4(
.number_in_stubinLink1(SL1_L4D4_VMR_L4D4_number),
.read_add_stubinLink1(SL1_L4D4_VMR_L4D4_read_add),
.stubinLink1(SL1_L4D4_VMR_L4D4),
.number_in_stubinLink2(SL2_L4D4_VMR_L4D4_number),
.read_add_stubinLink2(SL2_L4D4_VMR_L4D4_read_add),
.stubinLink2(SL2_L4D4_VMR_L4D4),
.number_in_stubinLink3(SL3_L4D4_VMR_L4D4_number),
.read_add_stubinLink3(SL3_L4D4_VMR_L4D4_read_add),
.stubinLink3(SL3_L4D4_VMR_L4D4),
.vmstuboutPHI1X1n1(VMR_L4D4_VMS_L4D4PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L4D4_VMS_L4D4PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L4D4_VMS_L4D4PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L4D4_VMS_L4D4PHI1X1n4),
.vmstuboutPHI2X1n1(VMR_L4D4_VMS_L4D4PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L4D4_VMS_L4D4PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L4D4_VMS_L4D4PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L4D4_VMS_L4D4PHI2X1n4),
.vmstuboutPHI2X1n5(VMR_L4D4_VMS_L4D4PHI2X1n5),
.vmstuboutPHI2X1n6(VMR_L4D4_VMS_L4D4PHI2X1n6),
.vmstuboutPHI3X1n1(VMR_L4D4_VMS_L4D4PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L4D4_VMS_L4D4PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L4D4_VMS_L4D4PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L4D4_VMS_L4D4PHI3X1n4),
.vmstuboutPHI3X1n5(VMR_L4D4_VMS_L4D4PHI3X1n5),
.vmstuboutPHI3X1n6(VMR_L4D4_VMS_L4D4PHI3X1n6),
.vmstuboutPHI4X1n1(VMR_L4D4_VMS_L4D4PHI4X1n1),
.vmstuboutPHI4X1n2(VMR_L4D4_VMS_L4D4PHI4X1n2),
.vmstuboutPHI4X1n3(VMR_L4D4_VMS_L4D4PHI4X1n3),
.vmstuboutPHI4X1n4(VMR_L4D4_VMS_L4D4PHI4X1n4),
.vmstuboutPHI1X2n1(VMR_L4D4_VMS_L4D4PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L4D4_VMS_L4D4PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L4D4_VMS_L4D4PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L4D4_VMS_L4D4PHI1X2n4),
.vmstuboutPHI2X2n1(VMR_L4D4_VMS_L4D4PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L4D4_VMS_L4D4PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L4D4_VMS_L4D4PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L4D4_VMS_L4D4PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L4D4_VMS_L4D4PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L4D4_VMS_L4D4PHI2X2n6),
.vmstuboutPHI3X2n1(VMR_L4D4_VMS_L4D4PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L4D4_VMS_L4D4PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L4D4_VMS_L4D4PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L4D4_VMS_L4D4PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L4D4_VMS_L4D4PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L4D4_VMS_L4D4PHI3X2n6),
.vmstuboutPHI4X2n1(VMR_L4D4_VMS_L4D4PHI4X2n1),
.vmstuboutPHI4X2n2(VMR_L4D4_VMS_L4D4PHI4X2n2),
.vmstuboutPHI4X2n3(VMR_L4D4_VMS_L4D4PHI4X2n3),
.vmstuboutPHI4X2n4(VMR_L4D4_VMS_L4D4PHI4X2n4),
.allstuboutn1(VMR_L4D4_AS_L4D4n1),
.allstuboutn2(VMR_L4D4_AS_L4D4n2),
.allstuboutn3(VMR_L4D4_AS_L4D4n3),
.allstuboutn4(VMR_L4D4_AS_L4D4n4),
.vmstuboutPHI1X1n1_wr_en(VMR_L4D4_VMS_L4D4PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L4D4_VMS_L4D4PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L4D4_VMS_L4D4PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L4D4_VMS_L4D4PHI1X1n4_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L4D4_VMS_L4D4PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L4D4_VMS_L4D4PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L4D4_VMS_L4D4PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L4D4_VMS_L4D4PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMR_L4D4_VMS_L4D4PHI2X1n5_wr_en),
.vmstuboutPHI2X1n6_wr_en(VMR_L4D4_VMS_L4D4PHI2X1n6_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L4D4_VMS_L4D4PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L4D4_VMS_L4D4PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L4D4_VMS_L4D4PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L4D4_VMS_L4D4PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMR_L4D4_VMS_L4D4PHI3X1n5_wr_en),
.vmstuboutPHI3X1n6_wr_en(VMR_L4D4_VMS_L4D4PHI3X1n6_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMR_L4D4_VMS_L4D4PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMR_L4D4_VMS_L4D4PHI4X1n2_wr_en),
.vmstuboutPHI4X1n3_wr_en(VMR_L4D4_VMS_L4D4PHI4X1n3_wr_en),
.vmstuboutPHI4X1n4_wr_en(VMR_L4D4_VMS_L4D4PHI4X1n4_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L4D4_VMS_L4D4PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L4D4_VMS_L4D4PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L4D4_VMS_L4D4PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L4D4_VMS_L4D4PHI1X2n4_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L4D4_VMS_L4D4PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L4D4_VMS_L4D4PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L4D4_VMS_L4D4PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L4D4_VMS_L4D4PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L4D4_VMS_L4D4PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L4D4_VMS_L4D4PHI2X2n6_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L4D4_VMS_L4D4PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L4D4_VMS_L4D4PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L4D4_VMS_L4D4PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L4D4_VMS_L4D4PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L4D4_VMS_L4D4PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L4D4_VMS_L4D4PHI3X2n6_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMR_L4D4_VMS_L4D4PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMR_L4D4_VMS_L4D4PHI4X2n2_wr_en),
.vmstuboutPHI4X2n3_wr_en(VMR_L4D4_VMS_L4D4PHI4X2n3_wr_en),
.vmstuboutPHI4X2n4_wr_en(VMR_L4D4_VMS_L4D4PHI4X2n4_wr_en),
.valid_data1(VMR_L4D4_AS_L4D4n1_wr_en),
.valid_data2(VMR_L4D4_AS_L4D4n2_wr_en),
.valid_data3(VMR_L4D4_AS_L4D4n3_wr_en),
.valid_data4(VMR_L4D4_AS_L4D4n4_wr_en),
.start(SL1_L4D4_start),
.done(VMR_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b0,1'b1) VMR_L5D3(
.number_in_stubinLink1(SL1_L5D3_VMR_L5D3_number),
.read_add_stubinLink1(SL1_L5D3_VMR_L5D3_read_add),
.stubinLink1(SL1_L5D3_VMR_L5D3),
.number_in_stubinLink2(SL2_L5D3_VMR_L5D3_number),
.read_add_stubinLink2(SL2_L5D3_VMR_L5D3_read_add),
.stubinLink2(SL2_L5D3_VMR_L5D3),
.number_in_stubinLink3(SL3_L5D3_VMR_L5D3_number),
.read_add_stubinLink3(SL3_L5D3_VMR_L5D3_read_add),
.stubinLink3(SL3_L5D3_VMR_L5D3),
.vmstuboutPHI1X1n1(VMR_L5D3_VMS_L5D3PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L5D3_VMS_L5D3PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L5D3_VMS_L5D3PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L5D3_VMS_L5D3PHI1X1n4),
.vmstuboutPHI1X1n5(VMR_L5D3_VMS_L5D3PHI1X1n5),
.vmstuboutPHI1X1n6(VMR_L5D3_VMS_L5D3PHI1X1n6),
.vmstuboutPHI2X1n1(VMR_L5D3_VMS_L5D3PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L5D3_VMS_L5D3PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L5D3_VMS_L5D3PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L5D3_VMS_L5D3PHI2X1n4),
.vmstuboutPHI2X1n5(VMR_L5D3_VMS_L5D3PHI2X1n5),
.vmstuboutPHI2X1n6(VMR_L5D3_VMS_L5D3PHI2X1n6),
.vmstuboutPHI3X1n1(VMR_L5D3_VMS_L5D3PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L5D3_VMS_L5D3PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L5D3_VMS_L5D3PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L5D3_VMS_L5D3PHI3X1n4),
.vmstuboutPHI3X1n5(VMR_L5D3_VMS_L5D3PHI3X1n5),
.vmstuboutPHI3X1n6(VMR_L5D3_VMS_L5D3PHI3X1n6),
.vmstuboutPHI1X2n1(VMR_L5D3_VMS_L5D3PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L5D3_VMS_L5D3PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L5D3_VMS_L5D3PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L5D3_VMS_L5D3PHI1X2n4),
.vmstuboutPHI1X2n5(VMR_L5D3_VMS_L5D3PHI1X2n5),
.vmstuboutPHI1X2n6(VMR_L5D3_VMS_L5D3PHI1X2n6),
.vmstuboutPHI2X2n1(VMR_L5D3_VMS_L5D3PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L5D3_VMS_L5D3PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L5D3_VMS_L5D3PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L5D3_VMS_L5D3PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L5D3_VMS_L5D3PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L5D3_VMS_L5D3PHI2X2n6),
.vmstuboutPHI3X2n1(VMR_L5D3_VMS_L5D3PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L5D3_VMS_L5D3PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L5D3_VMS_L5D3PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L5D3_VMS_L5D3PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L5D3_VMS_L5D3PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L5D3_VMS_L5D3PHI3X2n6),
.allstuboutn1(VMR_L5D3_AS_L5D3n1),
.allstuboutn2(VMR_L5D3_AS_L5D3n2),
.allstuboutn3(VMR_L5D3_AS_L5D3n3),
.allstuboutn4(VMR_L5D3_AS_L5D3n4),
.vmstuboutPHI1X1n1_wr_en(VMR_L5D3_VMS_L5D3PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L5D3_VMS_L5D3PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L5D3_VMS_L5D3PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L5D3_VMS_L5D3PHI1X1n4_wr_en),
.vmstuboutPHI1X1n5_wr_en(VMR_L5D3_VMS_L5D3PHI1X1n5_wr_en),
.vmstuboutPHI1X1n6_wr_en(VMR_L5D3_VMS_L5D3PHI1X1n6_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L5D3_VMS_L5D3PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L5D3_VMS_L5D3PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L5D3_VMS_L5D3PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L5D3_VMS_L5D3PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMR_L5D3_VMS_L5D3PHI2X1n5_wr_en),
.vmstuboutPHI2X1n6_wr_en(VMR_L5D3_VMS_L5D3PHI2X1n6_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L5D3_VMS_L5D3PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L5D3_VMS_L5D3PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L5D3_VMS_L5D3PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L5D3_VMS_L5D3PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMR_L5D3_VMS_L5D3PHI3X1n5_wr_en),
.vmstuboutPHI3X1n6_wr_en(VMR_L5D3_VMS_L5D3PHI3X1n6_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L5D3_VMS_L5D3PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L5D3_VMS_L5D3PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L5D3_VMS_L5D3PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L5D3_VMS_L5D3PHI1X2n4_wr_en),
.vmstuboutPHI1X2n5_wr_en(VMR_L5D3_VMS_L5D3PHI1X2n5_wr_en),
.vmstuboutPHI1X2n6_wr_en(VMR_L5D3_VMS_L5D3PHI1X2n6_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L5D3_VMS_L5D3PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L5D3_VMS_L5D3PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L5D3_VMS_L5D3PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L5D3_VMS_L5D3PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L5D3_VMS_L5D3PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L5D3_VMS_L5D3PHI2X2n6_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L5D3_VMS_L5D3PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L5D3_VMS_L5D3PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L5D3_VMS_L5D3PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L5D3_VMS_L5D3PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L5D3_VMS_L5D3PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L5D3_VMS_L5D3PHI3X2n6_wr_en),
.valid_data1(VMR_L5D3_AS_L5D3n1_wr_en),
.valid_data2(VMR_L5D3_AS_L5D3n2_wr_en),
.valid_data3(VMR_L5D3_AS_L5D3n3_wr_en),
.valid_data4(VMR_L5D3_AS_L5D3n4_wr_en),
.start(SL1_L5D3_start),
.done(VMR_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b0,1'b1) VMR_L5D4(
.number_in_stubinLink1(SL1_L5D4_VMR_L5D4_number),
.read_add_stubinLink1(SL1_L5D4_VMR_L5D4_read_add),
.stubinLink1(SL1_L5D4_VMR_L5D4),
.number_in_stubinLink2(SL2_L5D4_VMR_L5D4_number),
.read_add_stubinLink2(SL2_L5D4_VMR_L5D4_read_add),
.stubinLink2(SL2_L5D4_VMR_L5D4),
.number_in_stubinLink3(SL3_L5D4_VMR_L5D4_number),
.read_add_stubinLink3(SL3_L5D4_VMR_L5D4_read_add),
.stubinLink3(SL3_L5D4_VMR_L5D4),
.vmstuboutPHI1X1n1(VMR_L5D4_VMS_L5D4PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L5D4_VMS_L5D4PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L5D4_VMS_L5D4PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L5D4_VMS_L5D4PHI1X1n4),
.vmstuboutPHI1X1n5(VMR_L5D4_VMS_L5D4PHI1X1n5),
.vmstuboutPHI1X1n6(VMR_L5D4_VMS_L5D4PHI1X1n6),
.vmstuboutPHI2X1n1(VMR_L5D4_VMS_L5D4PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L5D4_VMS_L5D4PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L5D4_VMS_L5D4PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L5D4_VMS_L5D4PHI2X1n4),
.vmstuboutPHI2X1n5(VMR_L5D4_VMS_L5D4PHI2X1n5),
.vmstuboutPHI2X1n6(VMR_L5D4_VMS_L5D4PHI2X1n6),
.vmstuboutPHI3X1n1(VMR_L5D4_VMS_L5D4PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L5D4_VMS_L5D4PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L5D4_VMS_L5D4PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L5D4_VMS_L5D4PHI3X1n4),
.vmstuboutPHI3X1n5(VMR_L5D4_VMS_L5D4PHI3X1n5),
.vmstuboutPHI3X1n6(VMR_L5D4_VMS_L5D4PHI3X1n6),
.vmstuboutPHI1X2n1(VMR_L5D4_VMS_L5D4PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L5D4_VMS_L5D4PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L5D4_VMS_L5D4PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L5D4_VMS_L5D4PHI1X2n4),
.vmstuboutPHI2X2n1(VMR_L5D4_VMS_L5D4PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L5D4_VMS_L5D4PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L5D4_VMS_L5D4PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L5D4_VMS_L5D4PHI2X2n4),
.vmstuboutPHI3X2n1(VMR_L5D4_VMS_L5D4PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L5D4_VMS_L5D4PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L5D4_VMS_L5D4PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L5D4_VMS_L5D4PHI3X2n4),
.allstuboutn1(VMR_L5D4_AS_L5D4n1),
.allstuboutn2(VMR_L5D4_AS_L5D4n2),
.allstuboutn3(VMR_L5D4_AS_L5D4n3),
.vmstuboutPHI1X1n1_wr_en(VMR_L5D4_VMS_L5D4PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L5D4_VMS_L5D4PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L5D4_VMS_L5D4PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L5D4_VMS_L5D4PHI1X1n4_wr_en),
.vmstuboutPHI1X1n5_wr_en(VMR_L5D4_VMS_L5D4PHI1X1n5_wr_en),
.vmstuboutPHI1X1n6_wr_en(VMR_L5D4_VMS_L5D4PHI1X1n6_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L5D4_VMS_L5D4PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L5D4_VMS_L5D4PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L5D4_VMS_L5D4PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L5D4_VMS_L5D4PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMR_L5D4_VMS_L5D4PHI2X1n5_wr_en),
.vmstuboutPHI2X1n6_wr_en(VMR_L5D4_VMS_L5D4PHI2X1n6_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L5D4_VMS_L5D4PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L5D4_VMS_L5D4PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L5D4_VMS_L5D4PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L5D4_VMS_L5D4PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMR_L5D4_VMS_L5D4PHI3X1n5_wr_en),
.vmstuboutPHI3X1n6_wr_en(VMR_L5D4_VMS_L5D4PHI3X1n6_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L5D4_VMS_L5D4PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L5D4_VMS_L5D4PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L5D4_VMS_L5D4PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L5D4_VMS_L5D4PHI1X2n4_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L5D4_VMS_L5D4PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L5D4_VMS_L5D4PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L5D4_VMS_L5D4PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L5D4_VMS_L5D4PHI2X2n4_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L5D4_VMS_L5D4PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L5D4_VMS_L5D4PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L5D4_VMS_L5D4PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L5D4_VMS_L5D4PHI3X2n4_wr_en),
.valid_data1(VMR_L5D4_AS_L5D4n1_wr_en),
.valid_data2(VMR_L5D4_AS_L5D4n2_wr_en),
.valid_data3(VMR_L5D4_AS_L5D4n3_wr_en),
.start(SL1_L5D4_start),
.done(VMR_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b0,1'b0) VMR_L6D3(
.number_in_stubinLink1(SL1_L6D3_VMR_L6D3_number),
.read_add_stubinLink1(SL1_L6D3_VMR_L6D3_read_add),
.stubinLink1(SL1_L6D3_VMR_L6D3),
.number_in_stubinLink2(SL2_L6D3_VMR_L6D3_number),
.read_add_stubinLink2(SL2_L6D3_VMR_L6D3_read_add),
.stubinLink2(SL2_L6D3_VMR_L6D3),
.number_in_stubinLink3(SL3_L6D3_VMR_L6D3_number),
.read_add_stubinLink3(SL3_L6D3_VMR_L6D3_read_add),
.stubinLink3(SL3_L6D3_VMR_L6D3),
.vmstuboutPHI1X1n1(VMR_L6D3_VMS_L6D3PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L6D3_VMS_L6D3PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L6D3_VMS_L6D3PHI1X1n3),
.vmstuboutPHI2X1n1(VMR_L6D3_VMS_L6D3PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L6D3_VMS_L6D3PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L6D3_VMS_L6D3PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L6D3_VMS_L6D3PHI2X1n4),
.vmstuboutPHI3X1n1(VMR_L6D3_VMS_L6D3PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L6D3_VMS_L6D3PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L6D3_VMS_L6D3PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L6D3_VMS_L6D3PHI3X1n4),
.vmstuboutPHI4X1n1(VMR_L6D3_VMS_L6D3PHI4X1n1),
.vmstuboutPHI4X1n2(VMR_L6D3_VMS_L6D3PHI4X1n2),
.vmstuboutPHI4X1n3(VMR_L6D3_VMS_L6D3PHI4X1n3),
.vmstuboutPHI1X2n1(VMR_L6D3_VMS_L6D3PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L6D3_VMS_L6D3PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L6D3_VMS_L6D3PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L6D3_VMS_L6D3PHI1X2n4),
.vmstuboutPHI2X2n1(VMR_L6D3_VMS_L6D3PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L6D3_VMS_L6D3PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L6D3_VMS_L6D3PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L6D3_VMS_L6D3PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L6D3_VMS_L6D3PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L6D3_VMS_L6D3PHI2X2n6),
.vmstuboutPHI3X2n1(VMR_L6D3_VMS_L6D3PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L6D3_VMS_L6D3PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L6D3_VMS_L6D3PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L6D3_VMS_L6D3PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L6D3_VMS_L6D3PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L6D3_VMS_L6D3PHI3X2n6),
.vmstuboutPHI4X2n1(VMR_L6D3_VMS_L6D3PHI4X2n1),
.vmstuboutPHI4X2n2(VMR_L6D3_VMS_L6D3PHI4X2n2),
.vmstuboutPHI4X2n3(VMR_L6D3_VMS_L6D3PHI4X2n3),
.vmstuboutPHI4X2n4(VMR_L6D3_VMS_L6D3PHI4X2n4),
.allstuboutn1(VMR_L6D3_AS_L6D3n1),
.allstuboutn2(VMR_L6D3_AS_L6D3n2),
.allstuboutn3(VMR_L6D3_AS_L6D3n3),
.vmstuboutPHI1X1n1_wr_en(VMR_L6D3_VMS_L6D3PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L6D3_VMS_L6D3PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L6D3_VMS_L6D3PHI1X1n3_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L6D3_VMS_L6D3PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L6D3_VMS_L6D3PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L6D3_VMS_L6D3PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L6D3_VMS_L6D3PHI2X1n4_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L6D3_VMS_L6D3PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L6D3_VMS_L6D3PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L6D3_VMS_L6D3PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L6D3_VMS_L6D3PHI3X1n4_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMR_L6D3_VMS_L6D3PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMR_L6D3_VMS_L6D3PHI4X1n2_wr_en),
.vmstuboutPHI4X1n3_wr_en(VMR_L6D3_VMS_L6D3PHI4X1n3_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L6D3_VMS_L6D3PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L6D3_VMS_L6D3PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L6D3_VMS_L6D3PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L6D3_VMS_L6D3PHI1X2n4_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L6D3_VMS_L6D3PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L6D3_VMS_L6D3PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L6D3_VMS_L6D3PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L6D3_VMS_L6D3PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L6D3_VMS_L6D3PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L6D3_VMS_L6D3PHI2X2n6_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L6D3_VMS_L6D3PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L6D3_VMS_L6D3PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L6D3_VMS_L6D3PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L6D3_VMS_L6D3PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L6D3_VMS_L6D3PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L6D3_VMS_L6D3PHI3X2n6_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMR_L6D3_VMS_L6D3PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMR_L6D3_VMS_L6D3PHI4X2n2_wr_en),
.vmstuboutPHI4X2n3_wr_en(VMR_L6D3_VMS_L6D3PHI4X2n3_wr_en),
.vmstuboutPHI4X2n4_wr_en(VMR_L6D3_VMS_L6D3PHI4X2n4_wr_en),
.valid_data1(VMR_L6D3_AS_L6D3n1_wr_en),
.valid_data2(VMR_L6D3_AS_L6D3n2_wr_en),
.valid_data3(VMR_L6D3_AS_L6D3n3_wr_en),
.start(SL1_L6D3_start),
.done(VMR_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

VMRouter #(1'b0,1'b0) VMR_L6D4(
.number_in_stubinLink1(SL1_L6D4_VMR_L6D4_number),
.read_add_stubinLink1(SL1_L6D4_VMR_L6D4_read_add),
.stubinLink1(SL1_L6D4_VMR_L6D4),
.number_in_stubinLink2(SL2_L6D4_VMR_L6D4_number),
.read_add_stubinLink2(SL2_L6D4_VMR_L6D4_read_add),
.stubinLink2(SL2_L6D4_VMR_L6D4),
.number_in_stubinLink3(SL3_L6D4_VMR_L6D4_number),
.read_add_stubinLink3(SL3_L6D4_VMR_L6D4_read_add),
.stubinLink3(SL3_L6D4_VMR_L6D4),
.vmstuboutPHI1X1n1(VMR_L6D4_VMS_L6D4PHI1X1n1),
.vmstuboutPHI1X1n2(VMR_L6D4_VMS_L6D4PHI1X1n2),
.vmstuboutPHI1X1n3(VMR_L6D4_VMS_L6D4PHI1X1n3),
.vmstuboutPHI1X1n4(VMR_L6D4_VMS_L6D4PHI1X1n4),
.vmstuboutPHI2X1n1(VMR_L6D4_VMS_L6D4PHI2X1n1),
.vmstuboutPHI2X1n2(VMR_L6D4_VMS_L6D4PHI2X1n2),
.vmstuboutPHI2X1n3(VMR_L6D4_VMS_L6D4PHI2X1n3),
.vmstuboutPHI2X1n4(VMR_L6D4_VMS_L6D4PHI2X1n4),
.vmstuboutPHI2X1n5(VMR_L6D4_VMS_L6D4PHI2X1n5),
.vmstuboutPHI2X1n6(VMR_L6D4_VMS_L6D4PHI2X1n6),
.vmstuboutPHI3X1n1(VMR_L6D4_VMS_L6D4PHI3X1n1),
.vmstuboutPHI3X1n2(VMR_L6D4_VMS_L6D4PHI3X1n2),
.vmstuboutPHI3X1n3(VMR_L6D4_VMS_L6D4PHI3X1n3),
.vmstuboutPHI3X1n4(VMR_L6D4_VMS_L6D4PHI3X1n4),
.vmstuboutPHI3X1n5(VMR_L6D4_VMS_L6D4PHI3X1n5),
.vmstuboutPHI3X1n6(VMR_L6D4_VMS_L6D4PHI3X1n6),
.vmstuboutPHI4X1n1(VMR_L6D4_VMS_L6D4PHI4X1n1),
.vmstuboutPHI4X1n2(VMR_L6D4_VMS_L6D4PHI4X1n2),
.vmstuboutPHI4X1n3(VMR_L6D4_VMS_L6D4PHI4X1n3),
.vmstuboutPHI4X1n4(VMR_L6D4_VMS_L6D4PHI4X1n4),
.vmstuboutPHI1X2n1(VMR_L6D4_VMS_L6D4PHI1X2n1),
.vmstuboutPHI1X2n2(VMR_L6D4_VMS_L6D4PHI1X2n2),
.vmstuboutPHI1X2n3(VMR_L6D4_VMS_L6D4PHI1X2n3),
.vmstuboutPHI1X2n4(VMR_L6D4_VMS_L6D4PHI1X2n4),
.vmstuboutPHI2X2n1(VMR_L6D4_VMS_L6D4PHI2X2n1),
.vmstuboutPHI2X2n2(VMR_L6D4_VMS_L6D4PHI2X2n2),
.vmstuboutPHI2X2n3(VMR_L6D4_VMS_L6D4PHI2X2n3),
.vmstuboutPHI2X2n4(VMR_L6D4_VMS_L6D4PHI2X2n4),
.vmstuboutPHI2X2n5(VMR_L6D4_VMS_L6D4PHI2X2n5),
.vmstuboutPHI2X2n6(VMR_L6D4_VMS_L6D4PHI2X2n6),
.vmstuboutPHI3X2n1(VMR_L6D4_VMS_L6D4PHI3X2n1),
.vmstuboutPHI3X2n2(VMR_L6D4_VMS_L6D4PHI3X2n2),
.vmstuboutPHI3X2n3(VMR_L6D4_VMS_L6D4PHI3X2n3),
.vmstuboutPHI3X2n4(VMR_L6D4_VMS_L6D4PHI3X2n4),
.vmstuboutPHI3X2n5(VMR_L6D4_VMS_L6D4PHI3X2n5),
.vmstuboutPHI3X2n6(VMR_L6D4_VMS_L6D4PHI3X2n6),
.vmstuboutPHI4X2n1(VMR_L6D4_VMS_L6D4PHI4X2n1),
.vmstuboutPHI4X2n2(VMR_L6D4_VMS_L6D4PHI4X2n2),
.vmstuboutPHI4X2n3(VMR_L6D4_VMS_L6D4PHI4X2n3),
.vmstuboutPHI4X2n4(VMR_L6D4_VMS_L6D4PHI4X2n4),
.allstuboutn1(VMR_L6D4_AS_L6D4n1),
.allstuboutn2(VMR_L6D4_AS_L6D4n2),
.allstuboutn3(VMR_L6D4_AS_L6D4n3),
.allstuboutn4(VMR_L6D4_AS_L6D4n4),
.vmstuboutPHI1X1n1_wr_en(VMR_L6D4_VMS_L6D4PHI1X1n1_wr_en),
.vmstuboutPHI1X1n2_wr_en(VMR_L6D4_VMS_L6D4PHI1X1n2_wr_en),
.vmstuboutPHI1X1n3_wr_en(VMR_L6D4_VMS_L6D4PHI1X1n3_wr_en),
.vmstuboutPHI1X1n4_wr_en(VMR_L6D4_VMS_L6D4PHI1X1n4_wr_en),
.vmstuboutPHI2X1n1_wr_en(VMR_L6D4_VMS_L6D4PHI2X1n1_wr_en),
.vmstuboutPHI2X1n2_wr_en(VMR_L6D4_VMS_L6D4PHI2X1n2_wr_en),
.vmstuboutPHI2X1n3_wr_en(VMR_L6D4_VMS_L6D4PHI2X1n3_wr_en),
.vmstuboutPHI2X1n4_wr_en(VMR_L6D4_VMS_L6D4PHI2X1n4_wr_en),
.vmstuboutPHI2X1n5_wr_en(VMR_L6D4_VMS_L6D4PHI2X1n5_wr_en),
.vmstuboutPHI2X1n6_wr_en(VMR_L6D4_VMS_L6D4PHI2X1n6_wr_en),
.vmstuboutPHI3X1n1_wr_en(VMR_L6D4_VMS_L6D4PHI3X1n1_wr_en),
.vmstuboutPHI3X1n2_wr_en(VMR_L6D4_VMS_L6D4PHI3X1n2_wr_en),
.vmstuboutPHI3X1n3_wr_en(VMR_L6D4_VMS_L6D4PHI3X1n3_wr_en),
.vmstuboutPHI3X1n4_wr_en(VMR_L6D4_VMS_L6D4PHI3X1n4_wr_en),
.vmstuboutPHI3X1n5_wr_en(VMR_L6D4_VMS_L6D4PHI3X1n5_wr_en),
.vmstuboutPHI3X1n6_wr_en(VMR_L6D4_VMS_L6D4PHI3X1n6_wr_en),
.vmstuboutPHI4X1n1_wr_en(VMR_L6D4_VMS_L6D4PHI4X1n1_wr_en),
.vmstuboutPHI4X1n2_wr_en(VMR_L6D4_VMS_L6D4PHI4X1n2_wr_en),
.vmstuboutPHI4X1n3_wr_en(VMR_L6D4_VMS_L6D4PHI4X1n3_wr_en),
.vmstuboutPHI4X1n4_wr_en(VMR_L6D4_VMS_L6D4PHI4X1n4_wr_en),
.vmstuboutPHI1X2n1_wr_en(VMR_L6D4_VMS_L6D4PHI1X2n1_wr_en),
.vmstuboutPHI1X2n2_wr_en(VMR_L6D4_VMS_L6D4PHI1X2n2_wr_en),
.vmstuboutPHI1X2n3_wr_en(VMR_L6D4_VMS_L6D4PHI1X2n3_wr_en),
.vmstuboutPHI1X2n4_wr_en(VMR_L6D4_VMS_L6D4PHI1X2n4_wr_en),
.vmstuboutPHI2X2n1_wr_en(VMR_L6D4_VMS_L6D4PHI2X2n1_wr_en),
.vmstuboutPHI2X2n2_wr_en(VMR_L6D4_VMS_L6D4PHI2X2n2_wr_en),
.vmstuboutPHI2X2n3_wr_en(VMR_L6D4_VMS_L6D4PHI2X2n3_wr_en),
.vmstuboutPHI2X2n4_wr_en(VMR_L6D4_VMS_L6D4PHI2X2n4_wr_en),
.vmstuboutPHI2X2n5_wr_en(VMR_L6D4_VMS_L6D4PHI2X2n5_wr_en),
.vmstuboutPHI2X2n6_wr_en(VMR_L6D4_VMS_L6D4PHI2X2n6_wr_en),
.vmstuboutPHI3X2n1_wr_en(VMR_L6D4_VMS_L6D4PHI3X2n1_wr_en),
.vmstuboutPHI3X2n2_wr_en(VMR_L6D4_VMS_L6D4PHI3X2n2_wr_en),
.vmstuboutPHI3X2n3_wr_en(VMR_L6D4_VMS_L6D4PHI3X2n3_wr_en),
.vmstuboutPHI3X2n4_wr_en(VMR_L6D4_VMS_L6D4PHI3X2n4_wr_en),
.vmstuboutPHI3X2n5_wr_en(VMR_L6D4_VMS_L6D4PHI3X2n5_wr_en),
.vmstuboutPHI3X2n6_wr_en(VMR_L6D4_VMS_L6D4PHI3X2n6_wr_en),
.vmstuboutPHI4X2n1_wr_en(VMR_L6D4_VMS_L6D4PHI4X2n1_wr_en),
.vmstuboutPHI4X2n2_wr_en(VMR_L6D4_VMS_L6D4PHI4X2n2_wr_en),
.vmstuboutPHI4X2n3_wr_en(VMR_L6D4_VMS_L6D4PHI4X2n3_wr_en),
.vmstuboutPHI4X2n4_wr_en(VMR_L6D4_VMS_L6D4PHI4X2n4_wr_en),
.valid_data1(VMR_L6D4_AS_L6D4n1_wr_en),
.valid_data2(VMR_L6D4_AS_L6D4n2_wr_en),
.valid_data3(VMR_L6D4_AS_L6D4n3_wr_en),
.valid_data4(VMR_L6D4_AS_L6D4n4_wr_en),
.start(SL1_L6D4_start),
.done(VMR_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X1_L2D3PHI1X1_phi.txt","TETable_TE_L1D3PHI1X1_L2D3PHI1X1_z.txt") TE_L1D3PHI1X1_L2D3PHI1X1(
.number_in_innervmstubin(VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_number),
.read_add_innervmstubin(VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_read_add),
.innervmstubin(VMS_L1D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1),
.number_in_outervmstubin(VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_number),
.read_add_outervmstubin(VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1_read_add),
.outervmstubin(VMS_L2D3PHI1X1n1_TE_L1D3PHI1X1_L2D3PHI1X1),
.stubpairout(TE_L1D3PHI1X1_L2D3PHI1X1_SP_L1D3PHI1X1_L2D3PHI1X1),
.valid_data(TE_L1D3PHI1X1_L2D3PHI1X1_SP_L1D3PHI1X1_L2D3PHI1X1_wr_en),
.start(VMS_L1D3PHI1X1n1_start),
.done(TE_L1D3PHI1X1_L2D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X1_L2D3PHI2X1_phi.txt","TETable_TE_L1D3PHI1X1_L2D3PHI2X1_z.txt") TE_L1D3PHI1X1_L2D3PHI2X1(
.number_in_innervmstubin(VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1_number),
.read_add_innervmstubin(VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1_read_add),
.innervmstubin(VMS_L1D3PHI1X1n2_TE_L1D3PHI1X1_L2D3PHI2X1),
.number_in_outervmstubin(VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1_number),
.read_add_outervmstubin(VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1_read_add),
.outervmstubin(VMS_L2D3PHI2X1n1_TE_L1D3PHI1X1_L2D3PHI2X1),
.stubpairout(TE_L1D3PHI1X1_L2D3PHI2X1_SP_L1D3PHI1X1_L2D3PHI2X1),
.valid_data(TE_L1D3PHI1X1_L2D3PHI2X1_SP_L1D3PHI1X1_L2D3PHI2X1_wr_en),
.start(VMS_L1D3PHI1X1n2_start),
.done(TE_L1D3PHI1X1_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X1_L2D3PHI2X1_phi.txt","TETable_TE_L1D3PHI2X1_L2D3PHI2X1_z.txt") TE_L1D3PHI2X1_L2D3PHI2X1(
.number_in_outervmstubin(VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1_number),
.read_add_outervmstubin(VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1_read_add),
.outervmstubin(VMS_L2D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI2X1),
.number_in_innervmstubin(VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1_number),
.read_add_innervmstubin(VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1_read_add),
.innervmstubin(VMS_L1D3PHI2X1n1_TE_L1D3PHI2X1_L2D3PHI2X1),
.stubpairout(TE_L1D3PHI2X1_L2D3PHI2X1_SP_L1D3PHI2X1_L2D3PHI2X1),
.valid_data(TE_L1D3PHI2X1_L2D3PHI2X1_SP_L1D3PHI2X1_L2D3PHI2X1_wr_en),
.start(VMS_L2D3PHI2X1n2_start),
.done(TE_L1D3PHI2X1_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X1_L2D3PHI3X1_phi.txt","TETable_TE_L1D3PHI2X1_L2D3PHI3X1_z.txt") TE_L1D3PHI2X1_L2D3PHI3X1(
.number_in_innervmstubin(VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1_number),
.read_add_innervmstubin(VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1_read_add),
.innervmstubin(VMS_L1D3PHI2X1n2_TE_L1D3PHI2X1_L2D3PHI3X1),
.number_in_outervmstubin(VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1_number),
.read_add_outervmstubin(VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1_read_add),
.outervmstubin(VMS_L2D3PHI3X1n1_TE_L1D3PHI2X1_L2D3PHI3X1),
.stubpairout(TE_L1D3PHI2X1_L2D3PHI3X1_SP_L1D3PHI2X1_L2D3PHI3X1),
.valid_data(TE_L1D3PHI2X1_L2D3PHI3X1_SP_L1D3PHI2X1_L2D3PHI3X1_wr_en),
.start(VMS_L1D3PHI2X1n2_start),
.done(TE_L1D3PHI2X1_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X1_L2D3PHI3X1_phi.txt","TETable_TE_L1D3PHI3X1_L2D3PHI3X1_z.txt") TE_L1D3PHI3X1_L2D3PHI3X1(
.number_in_outervmstubin(VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1_number),
.read_add_outervmstubin(VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1_read_add),
.outervmstubin(VMS_L2D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI3X1),
.number_in_innervmstubin(VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1_number),
.read_add_innervmstubin(VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1_read_add),
.innervmstubin(VMS_L1D3PHI3X1n1_TE_L1D3PHI3X1_L2D3PHI3X1),
.stubpairout(TE_L1D3PHI3X1_L2D3PHI3X1_SP_L1D3PHI3X1_L2D3PHI3X1),
.valid_data(TE_L1D3PHI3X1_L2D3PHI3X1_SP_L1D3PHI3X1_L2D3PHI3X1_wr_en),
.start(VMS_L2D3PHI3X1n2_start),
.done(TE_L1D3PHI3X1_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X1_L2D3PHI4X1_phi.txt","TETable_TE_L1D3PHI3X1_L2D3PHI4X1_z.txt") TE_L1D3PHI3X1_L2D3PHI4X1(
.number_in_innervmstubin(VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1_number),
.read_add_innervmstubin(VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1_read_add),
.innervmstubin(VMS_L1D3PHI3X1n2_TE_L1D3PHI3X1_L2D3PHI4X1),
.number_in_outervmstubin(VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1_number),
.read_add_outervmstubin(VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1_read_add),
.outervmstubin(VMS_L2D3PHI4X1n1_TE_L1D3PHI3X1_L2D3PHI4X1),
.stubpairout(TE_L1D3PHI3X1_L2D3PHI4X1_SP_L1D3PHI3X1_L2D3PHI4X1),
.valid_data(TE_L1D3PHI3X1_L2D3PHI4X1_SP_L1D3PHI3X1_L2D3PHI4X1_wr_en),
.start(VMS_L1D3PHI3X1n2_start),
.done(TE_L1D3PHI3X1_L2D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X1_L2D3PHI1X2_phi.txt","TETable_TE_L1D3PHI1X1_L2D3PHI1X2_z.txt") TE_L1D3PHI1X1_L2D3PHI1X2(
.number_in_innervmstubin(VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2_number),
.read_add_innervmstubin(VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2_read_add),
.innervmstubin(VMS_L1D3PHI1X1n3_TE_L1D3PHI1X1_L2D3PHI1X2),
.number_in_outervmstubin(VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2_number),
.read_add_outervmstubin(VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2_read_add),
.outervmstubin(VMS_L2D3PHI1X2n1_TE_L1D3PHI1X1_L2D3PHI1X2),
.stubpairout(TE_L1D3PHI1X1_L2D3PHI1X2_SP_L1D3PHI1X1_L2D3PHI1X2),
.valid_data(TE_L1D3PHI1X1_L2D3PHI1X2_SP_L1D3PHI1X1_L2D3PHI1X2_wr_en),
.start(VMS_L1D3PHI1X1n3_start),
.done(TE_L1D3PHI1X1_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X1_L2D3PHI2X2_phi.txt","TETable_TE_L1D3PHI1X1_L2D3PHI2X2_z.txt") TE_L1D3PHI1X1_L2D3PHI2X2(
.number_in_innervmstubin(VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2_number),
.read_add_innervmstubin(VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2_read_add),
.innervmstubin(VMS_L1D3PHI1X1n4_TE_L1D3PHI1X1_L2D3PHI2X2),
.number_in_outervmstubin(VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2_number),
.read_add_outervmstubin(VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2_read_add),
.outervmstubin(VMS_L2D3PHI2X2n1_TE_L1D3PHI1X1_L2D3PHI2X2),
.stubpairout(TE_L1D3PHI1X1_L2D3PHI2X2_SP_L1D3PHI1X1_L2D3PHI2X2),
.valid_data(TE_L1D3PHI1X1_L2D3PHI2X2_SP_L1D3PHI1X1_L2D3PHI2X2_wr_en),
.start(VMS_L1D3PHI1X1n4_start),
.done(TE_L1D3PHI1X1_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X1_L2D3PHI2X2_phi.txt","TETable_TE_L1D3PHI2X1_L2D3PHI2X2_z.txt") TE_L1D3PHI2X1_L2D3PHI2X2(
.number_in_innervmstubin(VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2_number),
.read_add_innervmstubin(VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2_read_add),
.innervmstubin(VMS_L1D3PHI2X1n3_TE_L1D3PHI2X1_L2D3PHI2X2),
.number_in_outervmstubin(VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2_number),
.read_add_outervmstubin(VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2_read_add),
.outervmstubin(VMS_L2D3PHI2X2n2_TE_L1D3PHI2X1_L2D3PHI2X2),
.stubpairout(TE_L1D3PHI2X1_L2D3PHI2X2_SP_L1D3PHI2X1_L2D3PHI2X2),
.valid_data(TE_L1D3PHI2X1_L2D3PHI2X2_SP_L1D3PHI2X1_L2D3PHI2X2_wr_en),
.start(VMS_L1D3PHI2X1n3_start),
.done(TE_L1D3PHI2X1_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X1_L2D3PHI3X2_phi.txt","TETable_TE_L1D3PHI2X1_L2D3PHI3X2_z.txt") TE_L1D3PHI2X1_L2D3PHI3X2(
.number_in_innervmstubin(VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2_number),
.read_add_innervmstubin(VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2_read_add),
.innervmstubin(VMS_L1D3PHI2X1n4_TE_L1D3PHI2X1_L2D3PHI3X2),
.number_in_outervmstubin(VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2_number),
.read_add_outervmstubin(VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2_read_add),
.outervmstubin(VMS_L2D3PHI3X2n1_TE_L1D3PHI2X1_L2D3PHI3X2),
.stubpairout(TE_L1D3PHI2X1_L2D3PHI3X2_SP_L1D3PHI2X1_L2D3PHI3X2),
.valid_data(TE_L1D3PHI2X1_L2D3PHI3X2_SP_L1D3PHI2X1_L2D3PHI3X2_wr_en),
.start(VMS_L1D3PHI2X1n4_start),
.done(TE_L1D3PHI2X1_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X1_L2D3PHI3X2_phi.txt","TETable_TE_L1D3PHI3X1_L2D3PHI3X2_z.txt") TE_L1D3PHI3X1_L2D3PHI3X2(
.number_in_innervmstubin(VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2_number),
.read_add_innervmstubin(VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2_read_add),
.innervmstubin(VMS_L1D3PHI3X1n3_TE_L1D3PHI3X1_L2D3PHI3X2),
.number_in_outervmstubin(VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2_number),
.read_add_outervmstubin(VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2_read_add),
.outervmstubin(VMS_L2D3PHI3X2n2_TE_L1D3PHI3X1_L2D3PHI3X2),
.stubpairout(TE_L1D3PHI3X1_L2D3PHI3X2_SP_L1D3PHI3X1_L2D3PHI3X2),
.valid_data(TE_L1D3PHI3X1_L2D3PHI3X2_SP_L1D3PHI3X1_L2D3PHI3X2_wr_en),
.start(VMS_L1D3PHI3X1n3_start),
.done(TE_L1D3PHI3X1_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X1_L2D3PHI4X2_phi.txt","TETable_TE_L1D3PHI3X1_L2D3PHI4X2_z.txt") TE_L1D3PHI3X1_L2D3PHI4X2(
.number_in_innervmstubin(VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2_number),
.read_add_innervmstubin(VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2_read_add),
.innervmstubin(VMS_L1D3PHI3X1n4_TE_L1D3PHI3X1_L2D3PHI4X2),
.number_in_outervmstubin(VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2_number),
.read_add_outervmstubin(VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2_read_add),
.outervmstubin(VMS_L2D3PHI4X2n1_TE_L1D3PHI3X1_L2D3PHI4X2),
.stubpairout(TE_L1D3PHI3X1_L2D3PHI4X2_SP_L1D3PHI3X1_L2D3PHI4X2),
.valid_data(TE_L1D3PHI3X1_L2D3PHI4X2_SP_L1D3PHI3X1_L2D3PHI4X2_wr_en),
.start(VMS_L1D3PHI3X1n4_start),
.done(TE_L1D3PHI3X1_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X2_L2D3PHI1X2_phi.txt","TETable_TE_L1D3PHI1X2_L2D3PHI1X2_z.txt") TE_L1D3PHI1X2_L2D3PHI1X2(
.number_in_outervmstubin(VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2_number),
.read_add_outervmstubin(VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2_read_add),
.outervmstubin(VMS_L2D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI1X2),
.number_in_innervmstubin(VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2_number),
.read_add_innervmstubin(VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2_read_add),
.innervmstubin(VMS_L1D3PHI1X2n1_TE_L1D3PHI1X2_L2D3PHI1X2),
.stubpairout(TE_L1D3PHI1X2_L2D3PHI1X2_SP_L1D3PHI1X2_L2D3PHI1X2),
.valid_data(TE_L1D3PHI1X2_L2D3PHI1X2_SP_L1D3PHI1X2_L2D3PHI1X2_wr_en),
.start(VMS_L2D3PHI1X2n2_start),
.done(TE_L1D3PHI1X2_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X2_L2D3PHI2X2_phi.txt","TETable_TE_L1D3PHI1X2_L2D3PHI2X2_z.txt") TE_L1D3PHI1X2_L2D3PHI2X2(
.number_in_outervmstubin(VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2_number),
.read_add_outervmstubin(VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2_read_add),
.outervmstubin(VMS_L2D3PHI2X2n3_TE_L1D3PHI1X2_L2D3PHI2X2),
.number_in_innervmstubin(VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2_number),
.read_add_innervmstubin(VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2_read_add),
.innervmstubin(VMS_L1D3PHI1X2n2_TE_L1D3PHI1X2_L2D3PHI2X2),
.stubpairout(TE_L1D3PHI1X2_L2D3PHI2X2_SP_L1D3PHI1X2_L2D3PHI2X2),
.valid_data(TE_L1D3PHI1X2_L2D3PHI2X2_SP_L1D3PHI1X2_L2D3PHI2X2_wr_en),
.start(VMS_L2D3PHI2X2n3_start),
.done(TE_L1D3PHI1X2_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X2_L2D3PHI2X2_phi.txt","TETable_TE_L1D3PHI2X2_L2D3PHI2X2_z.txt") TE_L1D3PHI2X2_L2D3PHI2X2(
.number_in_outervmstubin(VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2_number),
.read_add_outervmstubin(VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2_read_add),
.outervmstubin(VMS_L2D3PHI2X2n4_TE_L1D3PHI2X2_L2D3PHI2X2),
.number_in_innervmstubin(VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2_number),
.read_add_innervmstubin(VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2_read_add),
.innervmstubin(VMS_L1D3PHI2X2n1_TE_L1D3PHI2X2_L2D3PHI2X2),
.stubpairout(TE_L1D3PHI2X2_L2D3PHI2X2_SP_L1D3PHI2X2_L2D3PHI2X2),
.valid_data(TE_L1D3PHI2X2_L2D3PHI2X2_SP_L1D3PHI2X2_L2D3PHI2X2_wr_en),
.start(VMS_L2D3PHI2X2n4_start),
.done(TE_L1D3PHI2X2_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X2_L2D3PHI3X2_phi.txt","TETable_TE_L1D3PHI2X2_L2D3PHI3X2_z.txt") TE_L1D3PHI2X2_L2D3PHI3X2(
.number_in_outervmstubin(VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2_number),
.read_add_outervmstubin(VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2_read_add),
.outervmstubin(VMS_L2D3PHI3X2n3_TE_L1D3PHI2X2_L2D3PHI3X2),
.number_in_innervmstubin(VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2_number),
.read_add_innervmstubin(VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2_read_add),
.innervmstubin(VMS_L1D3PHI2X2n2_TE_L1D3PHI2X2_L2D3PHI3X2),
.stubpairout(TE_L1D3PHI2X2_L2D3PHI3X2_SP_L1D3PHI2X2_L2D3PHI3X2),
.valid_data(TE_L1D3PHI2X2_L2D3PHI3X2_SP_L1D3PHI2X2_L2D3PHI3X2_wr_en),
.start(VMS_L2D3PHI3X2n3_start),
.done(TE_L1D3PHI2X2_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X2_L2D3PHI3X2_phi.txt","TETable_TE_L1D3PHI3X2_L2D3PHI3X2_z.txt") TE_L1D3PHI3X2_L2D3PHI3X2(
.number_in_outervmstubin(VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2_number),
.read_add_outervmstubin(VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2_read_add),
.outervmstubin(VMS_L2D3PHI3X2n4_TE_L1D3PHI3X2_L2D3PHI3X2),
.number_in_innervmstubin(VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2_number),
.read_add_innervmstubin(VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2_read_add),
.innervmstubin(VMS_L1D3PHI3X2n1_TE_L1D3PHI3X2_L2D3PHI3X2),
.stubpairout(TE_L1D3PHI3X2_L2D3PHI3X2_SP_L1D3PHI3X2_L2D3PHI3X2),
.valid_data(TE_L1D3PHI3X2_L2D3PHI3X2_SP_L1D3PHI3X2_L2D3PHI3X2_wr_en),
.start(VMS_L2D3PHI3X2n4_start),
.done(TE_L1D3PHI3X2_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X2_L2D3PHI4X2_phi.txt","TETable_TE_L1D3PHI3X2_L2D3PHI4X2_z.txt") TE_L1D3PHI3X2_L2D3PHI4X2(
.number_in_outervmstubin(VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_number),
.read_add_outervmstubin(VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_read_add),
.outervmstubin(VMS_L2D3PHI4X2n2_TE_L1D3PHI3X2_L2D3PHI4X2),
.number_in_innervmstubin(VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_number),
.read_add_innervmstubin(VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2_read_add),
.innervmstubin(VMS_L1D3PHI3X2n2_TE_L1D3PHI3X2_L2D3PHI4X2),
.stubpairout(TE_L1D3PHI3X2_L2D3PHI4X2_SP_L1D3PHI3X2_L2D3PHI4X2),
.valid_data(TE_L1D3PHI3X2_L2D3PHI4X2_SP_L1D3PHI3X2_L2D3PHI4X2_wr_en),
.start(VMS_L2D3PHI4X2n2_start),
.done(TE_L1D3PHI3X2_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X1_L2D4PHI1X1_phi.txt","TETable_TE_L1D3PHI1X1_L2D4PHI1X1_z.txt") TE_L1D3PHI1X1_L2D4PHI1X1(
.number_in_innervmstubin(VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1_number),
.read_add_innervmstubin(VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1_read_add),
.innervmstubin(VMS_L1D3PHI1X1n5_TE_L1D3PHI1X1_L2D4PHI1X1),
.number_in_outervmstubin(VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1_number),
.read_add_outervmstubin(VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1_read_add),
.outervmstubin(VMS_L2D4PHI1X1n1_TE_L1D3PHI1X1_L2D4PHI1X1),
.stubpairout(TE_L1D3PHI1X1_L2D4PHI1X1_SP_L1D3PHI1X1_L2D4PHI1X1),
.valid_data(TE_L1D3PHI1X1_L2D4PHI1X1_SP_L1D3PHI1X1_L2D4PHI1X1_wr_en),
.start(VMS_L1D3PHI1X1n5_start),
.done(TE_L1D3PHI1X1_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X1_L2D4PHI2X1_phi.txt","TETable_TE_L1D3PHI1X1_L2D4PHI2X1_z.txt") TE_L1D3PHI1X1_L2D4PHI2X1(
.number_in_innervmstubin(VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1_number),
.read_add_innervmstubin(VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1_read_add),
.innervmstubin(VMS_L1D3PHI1X1n6_TE_L1D3PHI1X1_L2D4PHI2X1),
.number_in_outervmstubin(VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1_number),
.read_add_outervmstubin(VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1_read_add),
.outervmstubin(VMS_L2D4PHI2X1n1_TE_L1D3PHI1X1_L2D4PHI2X1),
.stubpairout(TE_L1D3PHI1X1_L2D4PHI2X1_SP_L1D3PHI1X1_L2D4PHI2X1),
.valid_data(TE_L1D3PHI1X1_L2D4PHI2X1_SP_L1D3PHI1X1_L2D4PHI2X1_wr_en),
.start(VMS_L1D3PHI1X1n6_start),
.done(TE_L1D3PHI1X1_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X1_L2D4PHI2X1_phi.txt","TETable_TE_L1D3PHI2X1_L2D4PHI2X1_z.txt") TE_L1D3PHI2X1_L2D4PHI2X1(
.number_in_innervmstubin(VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1_number),
.read_add_innervmstubin(VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1_read_add),
.innervmstubin(VMS_L1D3PHI2X1n5_TE_L1D3PHI2X1_L2D4PHI2X1),
.number_in_outervmstubin(VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1_number),
.read_add_outervmstubin(VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1_read_add),
.outervmstubin(VMS_L2D4PHI2X1n2_TE_L1D3PHI2X1_L2D4PHI2X1),
.stubpairout(TE_L1D3PHI2X1_L2D4PHI2X1_SP_L1D3PHI2X1_L2D4PHI2X1),
.valid_data(TE_L1D3PHI2X1_L2D4PHI2X1_SP_L1D3PHI2X1_L2D4PHI2X1_wr_en),
.start(VMS_L1D3PHI2X1n5_start),
.done(TE_L1D3PHI2X1_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X1_L2D4PHI3X1_phi.txt","TETable_TE_L1D3PHI2X1_L2D4PHI3X1_z.txt") TE_L1D3PHI2X1_L2D4PHI3X1(
.number_in_innervmstubin(VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1_number),
.read_add_innervmstubin(VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1_read_add),
.innervmstubin(VMS_L1D3PHI2X1n6_TE_L1D3PHI2X1_L2D4PHI3X1),
.number_in_outervmstubin(VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1_number),
.read_add_outervmstubin(VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1_read_add),
.outervmstubin(VMS_L2D4PHI3X1n1_TE_L1D3PHI2X1_L2D4PHI3X1),
.stubpairout(TE_L1D3PHI2X1_L2D4PHI3X1_SP_L1D3PHI2X1_L2D4PHI3X1),
.valid_data(TE_L1D3PHI2X1_L2D4PHI3X1_SP_L1D3PHI2X1_L2D4PHI3X1_wr_en),
.start(VMS_L1D3PHI2X1n6_start),
.done(TE_L1D3PHI2X1_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X1_L2D4PHI3X1_phi.txt","TETable_TE_L1D3PHI3X1_L2D4PHI3X1_z.txt") TE_L1D3PHI3X1_L2D4PHI3X1(
.number_in_innervmstubin(VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1_number),
.read_add_innervmstubin(VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1_read_add),
.innervmstubin(VMS_L1D3PHI3X1n5_TE_L1D3PHI3X1_L2D4PHI3X1),
.number_in_outervmstubin(VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1_number),
.read_add_outervmstubin(VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1_read_add),
.outervmstubin(VMS_L2D4PHI3X1n2_TE_L1D3PHI3X1_L2D4PHI3X1),
.stubpairout(TE_L1D3PHI3X1_L2D4PHI3X1_SP_L1D3PHI3X1_L2D4PHI3X1),
.valid_data(TE_L1D3PHI3X1_L2D4PHI3X1_SP_L1D3PHI3X1_L2D4PHI3X1_wr_en),
.start(VMS_L1D3PHI3X1n5_start),
.done(TE_L1D3PHI3X1_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X1_L2D4PHI4X1_phi.txt","TETable_TE_L1D3PHI3X1_L2D4PHI4X1_z.txt") TE_L1D3PHI3X1_L2D4PHI4X1(
.number_in_innervmstubin(VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1_number),
.read_add_innervmstubin(VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1_read_add),
.innervmstubin(VMS_L1D3PHI3X1n6_TE_L1D3PHI3X1_L2D4PHI4X1),
.number_in_outervmstubin(VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1_number),
.read_add_outervmstubin(VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1_read_add),
.outervmstubin(VMS_L2D4PHI4X1n1_TE_L1D3PHI3X1_L2D4PHI4X1),
.stubpairout(TE_L1D3PHI3X1_L2D4PHI4X1_SP_L1D3PHI3X1_L2D4PHI4X1),
.valid_data(TE_L1D3PHI3X1_L2D4PHI4X1_SP_L1D3PHI3X1_L2D4PHI4X1_wr_en),
.start(VMS_L1D3PHI3X1n6_start),
.done(TE_L1D3PHI3X1_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X2_L2D4PHI1X1_phi.txt","TETable_TE_L1D3PHI1X2_L2D4PHI1X1_z.txt") TE_L1D3PHI1X2_L2D4PHI1X1(
.number_in_innervmstubin(VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1_number),
.read_add_innervmstubin(VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1_read_add),
.innervmstubin(VMS_L1D3PHI1X2n3_TE_L1D3PHI1X2_L2D4PHI1X1),
.number_in_outervmstubin(VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1_number),
.read_add_outervmstubin(VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1_read_add),
.outervmstubin(VMS_L2D4PHI1X1n2_TE_L1D3PHI1X2_L2D4PHI1X1),
.stubpairout(TE_L1D3PHI1X2_L2D4PHI1X1_SP_L1D3PHI1X2_L2D4PHI1X1),
.valid_data(TE_L1D3PHI1X2_L2D4PHI1X1_SP_L1D3PHI1X2_L2D4PHI1X1_wr_en),
.start(VMS_L1D3PHI1X2n3_start),
.done(TE_L1D3PHI1X2_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X2_L2D4PHI2X1_phi.txt","TETable_TE_L1D3PHI1X2_L2D4PHI2X1_z.txt") TE_L1D3PHI1X2_L2D4PHI2X1(
.number_in_innervmstubin(VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1_number),
.read_add_innervmstubin(VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1_read_add),
.innervmstubin(VMS_L1D3PHI1X2n4_TE_L1D3PHI1X2_L2D4PHI2X1),
.number_in_outervmstubin(VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1_number),
.read_add_outervmstubin(VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1_read_add),
.outervmstubin(VMS_L2D4PHI2X1n3_TE_L1D3PHI1X2_L2D4PHI2X1),
.stubpairout(TE_L1D3PHI1X2_L2D4PHI2X1_SP_L1D3PHI1X2_L2D4PHI2X1),
.valid_data(TE_L1D3PHI1X2_L2D4PHI2X1_SP_L1D3PHI1X2_L2D4PHI2X1_wr_en),
.start(VMS_L1D3PHI1X2n4_start),
.done(TE_L1D3PHI1X2_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X2_L2D4PHI2X1_phi.txt","TETable_TE_L1D3PHI2X2_L2D4PHI2X1_z.txt") TE_L1D3PHI2X2_L2D4PHI2X1(
.number_in_innervmstubin(VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1_number),
.read_add_innervmstubin(VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1_read_add),
.innervmstubin(VMS_L1D3PHI2X2n3_TE_L1D3PHI2X2_L2D4PHI2X1),
.number_in_outervmstubin(VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1_number),
.read_add_outervmstubin(VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1_read_add),
.outervmstubin(VMS_L2D4PHI2X1n4_TE_L1D3PHI2X2_L2D4PHI2X1),
.stubpairout(TE_L1D3PHI2X2_L2D4PHI2X1_SP_L1D3PHI2X2_L2D4PHI2X1),
.valid_data(TE_L1D3PHI2X2_L2D4PHI2X1_SP_L1D3PHI2X2_L2D4PHI2X1_wr_en),
.start(VMS_L1D3PHI2X2n3_start),
.done(TE_L1D3PHI2X2_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X2_L2D4PHI3X1_phi.txt","TETable_TE_L1D3PHI2X2_L2D4PHI3X1_z.txt") TE_L1D3PHI2X2_L2D4PHI3X1(
.number_in_innervmstubin(VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1_number),
.read_add_innervmstubin(VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1_read_add),
.innervmstubin(VMS_L1D3PHI2X2n4_TE_L1D3PHI2X2_L2D4PHI3X1),
.number_in_outervmstubin(VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1_number),
.read_add_outervmstubin(VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1_read_add),
.outervmstubin(VMS_L2D4PHI3X1n3_TE_L1D3PHI2X2_L2D4PHI3X1),
.stubpairout(TE_L1D3PHI2X2_L2D4PHI3X1_SP_L1D3PHI2X2_L2D4PHI3X1),
.valid_data(TE_L1D3PHI2X2_L2D4PHI3X1_SP_L1D3PHI2X2_L2D4PHI3X1_wr_en),
.start(VMS_L1D3PHI2X2n4_start),
.done(TE_L1D3PHI2X2_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X2_L2D4PHI3X1_phi.txt","TETable_TE_L1D3PHI3X2_L2D4PHI3X1_z.txt") TE_L1D3PHI3X2_L2D4PHI3X1(
.number_in_innervmstubin(VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1_number),
.read_add_innervmstubin(VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1_read_add),
.innervmstubin(VMS_L1D3PHI3X2n3_TE_L1D3PHI3X2_L2D4PHI3X1),
.number_in_outervmstubin(VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1_number),
.read_add_outervmstubin(VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1_read_add),
.outervmstubin(VMS_L2D4PHI3X1n4_TE_L1D3PHI3X2_L2D4PHI3X1),
.stubpairout(TE_L1D3PHI3X2_L2D4PHI3X1_SP_L1D3PHI3X2_L2D4PHI3X1),
.valid_data(TE_L1D3PHI3X2_L2D4PHI3X1_SP_L1D3PHI3X2_L2D4PHI3X1_wr_en),
.start(VMS_L1D3PHI3X2n3_start),
.done(TE_L1D3PHI3X2_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X2_L2D4PHI4X1_phi.txt","TETable_TE_L1D3PHI3X2_L2D4PHI4X1_z.txt") TE_L1D3PHI3X2_L2D4PHI4X1(
.number_in_innervmstubin(VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1_number),
.read_add_innervmstubin(VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1_read_add),
.innervmstubin(VMS_L1D3PHI3X2n4_TE_L1D3PHI3X2_L2D4PHI4X1),
.number_in_outervmstubin(VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1_number),
.read_add_outervmstubin(VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1_read_add),
.outervmstubin(VMS_L2D4PHI4X1n2_TE_L1D3PHI3X2_L2D4PHI4X1),
.stubpairout(TE_L1D3PHI3X2_L2D4PHI4X1_SP_L1D3PHI3X2_L2D4PHI4X1),
.valid_data(TE_L1D3PHI3X2_L2D4PHI4X1_SP_L1D3PHI3X2_L2D4PHI4X1_wr_en),
.start(VMS_L1D3PHI3X2n4_start),
.done(TE_L1D3PHI3X2_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X2_L2D4PHI1X2_phi.txt","TETable_TE_L1D3PHI1X2_L2D4PHI1X2_z.txt") TE_L1D3PHI1X2_L2D4PHI1X2(
.number_in_innervmstubin(VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2_number),
.read_add_innervmstubin(VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2_read_add),
.innervmstubin(VMS_L1D3PHI1X2n5_TE_L1D3PHI1X2_L2D4PHI1X2),
.number_in_outervmstubin(VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2_number),
.read_add_outervmstubin(VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2_read_add),
.outervmstubin(VMS_L2D4PHI1X2n1_TE_L1D3PHI1X2_L2D4PHI1X2),
.stubpairout(TE_L1D3PHI1X2_L2D4PHI1X2_SP_L1D3PHI1X2_L2D4PHI1X2),
.valid_data(TE_L1D3PHI1X2_L2D4PHI1X2_SP_L1D3PHI1X2_L2D4PHI1X2_wr_en),
.start(VMS_L1D3PHI1X2n5_start),
.done(TE_L1D3PHI1X2_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI1X2_L2D4PHI2X2_phi.txt","TETable_TE_L1D3PHI1X2_L2D4PHI2X2_z.txt") TE_L1D3PHI1X2_L2D4PHI2X2(
.number_in_innervmstubin(VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2_number),
.read_add_innervmstubin(VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2_read_add),
.innervmstubin(VMS_L1D3PHI1X2n6_TE_L1D3PHI1X2_L2D4PHI2X2),
.number_in_outervmstubin(VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2_number),
.read_add_outervmstubin(VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2_read_add),
.outervmstubin(VMS_L2D4PHI2X2n1_TE_L1D3PHI1X2_L2D4PHI2X2),
.stubpairout(TE_L1D3PHI1X2_L2D4PHI2X2_SP_L1D3PHI1X2_L2D4PHI2X2),
.valid_data(TE_L1D3PHI1X2_L2D4PHI2X2_SP_L1D3PHI1X2_L2D4PHI2X2_wr_en),
.start(VMS_L1D3PHI1X2n6_start),
.done(TE_L1D3PHI1X2_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X2_L2D4PHI2X2_phi.txt","TETable_TE_L1D3PHI2X2_L2D4PHI2X2_z.txt") TE_L1D3PHI2X2_L2D4PHI2X2(
.number_in_innervmstubin(VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2_number),
.read_add_innervmstubin(VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2_read_add),
.innervmstubin(VMS_L1D3PHI2X2n5_TE_L1D3PHI2X2_L2D4PHI2X2),
.number_in_outervmstubin(VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2_number),
.read_add_outervmstubin(VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2_read_add),
.outervmstubin(VMS_L2D4PHI2X2n2_TE_L1D3PHI2X2_L2D4PHI2X2),
.stubpairout(TE_L1D3PHI2X2_L2D4PHI2X2_SP_L1D3PHI2X2_L2D4PHI2X2),
.valid_data(TE_L1D3PHI2X2_L2D4PHI2X2_SP_L1D3PHI2X2_L2D4PHI2X2_wr_en),
.start(VMS_L1D3PHI2X2n5_start),
.done(TE_L1D3PHI2X2_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI2X2_L2D4PHI3X2_phi.txt","TETable_TE_L1D3PHI2X2_L2D4PHI3X2_z.txt") TE_L1D3PHI2X2_L2D4PHI3X2(
.number_in_innervmstubin(VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2_number),
.read_add_innervmstubin(VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2_read_add),
.innervmstubin(VMS_L1D3PHI2X2n6_TE_L1D3PHI2X2_L2D4PHI3X2),
.number_in_outervmstubin(VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2_number),
.read_add_outervmstubin(VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2_read_add),
.outervmstubin(VMS_L2D4PHI3X2n1_TE_L1D3PHI2X2_L2D4PHI3X2),
.stubpairout(TE_L1D3PHI2X2_L2D4PHI3X2_SP_L1D3PHI2X2_L2D4PHI3X2),
.valid_data(TE_L1D3PHI2X2_L2D4PHI3X2_SP_L1D3PHI2X2_L2D4PHI3X2_wr_en),
.start(VMS_L1D3PHI2X2n6_start),
.done(TE_L1D3PHI2X2_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X2_L2D4PHI3X2_phi.txt","TETable_TE_L1D3PHI3X2_L2D4PHI3X2_z.txt") TE_L1D3PHI3X2_L2D4PHI3X2(
.number_in_innervmstubin(VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2_number),
.read_add_innervmstubin(VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2_read_add),
.innervmstubin(VMS_L1D3PHI3X2n5_TE_L1D3PHI3X2_L2D4PHI3X2),
.number_in_outervmstubin(VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2_number),
.read_add_outervmstubin(VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2_read_add),
.outervmstubin(VMS_L2D4PHI3X2n2_TE_L1D3PHI3X2_L2D4PHI3X2),
.stubpairout(TE_L1D3PHI3X2_L2D4PHI3X2_SP_L1D3PHI3X2_L2D4PHI3X2),
.valid_data(TE_L1D3PHI3X2_L2D4PHI3X2_SP_L1D3PHI3X2_L2D4PHI3X2_wr_en),
.start(VMS_L1D3PHI3X2n5_start),
.done(TE_L1D3PHI3X2_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D3PHI3X2_L2D4PHI4X2_phi.txt","TETable_TE_L1D3PHI3X2_L2D4PHI4X2_z.txt") TE_L1D3PHI3X2_L2D4PHI4X2(
.number_in_innervmstubin(VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2_number),
.read_add_innervmstubin(VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2_read_add),
.innervmstubin(VMS_L1D3PHI3X2n6_TE_L1D3PHI3X2_L2D4PHI4X2),
.number_in_outervmstubin(VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2_number),
.read_add_outervmstubin(VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2_read_add),
.outervmstubin(VMS_L2D4PHI4X2n1_TE_L1D3PHI3X2_L2D4PHI4X2),
.stubpairout(TE_L1D3PHI3X2_L2D4PHI4X2_SP_L1D3PHI3X2_L2D4PHI4X2),
.valid_data(TE_L1D3PHI3X2_L2D4PHI4X2_SP_L1D3PHI3X2_L2D4PHI4X2_wr_en),
.start(VMS_L1D3PHI3X2n6_start),
.done(TE_L1D3PHI3X2_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D4PHI1X1_L2D4PHI1X2_phi.txt","TETable_TE_L1D4PHI1X1_L2D4PHI1X2_z.txt") TE_L1D4PHI1X1_L2D4PHI1X2(
.number_in_outervmstubin(VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2_number),
.read_add_outervmstubin(VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2_read_add),
.outervmstubin(VMS_L2D4PHI1X2n2_TE_L1D4PHI1X1_L2D4PHI1X2),
.number_in_innervmstubin(VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2_number),
.read_add_innervmstubin(VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2_read_add),
.innervmstubin(VMS_L1D4PHI1X1n1_TE_L1D4PHI1X1_L2D4PHI1X2),
.stubpairout(TE_L1D4PHI1X1_L2D4PHI1X2_SP_L1D4PHI1X1_L2D4PHI1X2),
.valid_data(TE_L1D4PHI1X1_L2D4PHI1X2_SP_L1D4PHI1X1_L2D4PHI1X2_wr_en),
.start(VMS_L2D4PHI1X2n2_start),
.done(TE_L1D4PHI1X1_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D4PHI1X1_L2D4PHI2X2_phi.txt","TETable_TE_L1D4PHI1X1_L2D4PHI2X2_z.txt") TE_L1D4PHI1X1_L2D4PHI2X2(
.number_in_outervmstubin(VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2_number),
.read_add_outervmstubin(VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2_read_add),
.outervmstubin(VMS_L2D4PHI2X2n3_TE_L1D4PHI1X1_L2D4PHI2X2),
.number_in_innervmstubin(VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2_number),
.read_add_innervmstubin(VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2_read_add),
.innervmstubin(VMS_L1D4PHI1X1n2_TE_L1D4PHI1X1_L2D4PHI2X2),
.stubpairout(TE_L1D4PHI1X1_L2D4PHI2X2_SP_L1D4PHI1X1_L2D4PHI2X2),
.valid_data(TE_L1D4PHI1X1_L2D4PHI2X2_SP_L1D4PHI1X1_L2D4PHI2X2_wr_en),
.start(VMS_L2D4PHI2X2n3_start),
.done(TE_L1D4PHI1X1_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D4PHI2X1_L2D4PHI2X2_phi.txt","TETable_TE_L1D4PHI2X1_L2D4PHI2X2_z.txt") TE_L1D4PHI2X1_L2D4PHI2X2(
.number_in_outervmstubin(VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2_number),
.read_add_outervmstubin(VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2_read_add),
.outervmstubin(VMS_L2D4PHI2X2n4_TE_L1D4PHI2X1_L2D4PHI2X2),
.number_in_innervmstubin(VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2_number),
.read_add_innervmstubin(VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2_read_add),
.innervmstubin(VMS_L1D4PHI2X1n1_TE_L1D4PHI2X1_L2D4PHI2X2),
.stubpairout(TE_L1D4PHI2X1_L2D4PHI2X2_SP_L1D4PHI2X1_L2D4PHI2X2),
.valid_data(TE_L1D4PHI2X1_L2D4PHI2X2_SP_L1D4PHI2X1_L2D4PHI2X2_wr_en),
.start(VMS_L2D4PHI2X2n4_start),
.done(TE_L1D4PHI2X1_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D4PHI2X1_L2D4PHI3X2_phi.txt","TETable_TE_L1D4PHI2X1_L2D4PHI3X2_z.txt") TE_L1D4PHI2X1_L2D4PHI3X2(
.number_in_outervmstubin(VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2_number),
.read_add_outervmstubin(VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2_read_add),
.outervmstubin(VMS_L2D4PHI3X2n3_TE_L1D4PHI2X1_L2D4PHI3X2),
.number_in_innervmstubin(VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2_number),
.read_add_innervmstubin(VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2_read_add),
.innervmstubin(VMS_L1D4PHI2X1n2_TE_L1D4PHI2X1_L2D4PHI3X2),
.stubpairout(TE_L1D4PHI2X1_L2D4PHI3X2_SP_L1D4PHI2X1_L2D4PHI3X2),
.valid_data(TE_L1D4PHI2X1_L2D4PHI3X2_SP_L1D4PHI2X1_L2D4PHI3X2_wr_en),
.start(VMS_L2D4PHI3X2n3_start),
.done(TE_L1D4PHI2X1_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D4PHI3X1_L2D4PHI3X2_phi.txt","TETable_TE_L1D4PHI3X1_L2D4PHI3X2_z.txt") TE_L1D4PHI3X1_L2D4PHI3X2(
.number_in_outervmstubin(VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2_number),
.read_add_outervmstubin(VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2_read_add),
.outervmstubin(VMS_L2D4PHI3X2n4_TE_L1D4PHI3X1_L2D4PHI3X2),
.number_in_innervmstubin(VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2_number),
.read_add_innervmstubin(VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2_read_add),
.innervmstubin(VMS_L1D4PHI3X1n1_TE_L1D4PHI3X1_L2D4PHI3X2),
.stubpairout(TE_L1D4PHI3X1_L2D4PHI3X2_SP_L1D4PHI3X1_L2D4PHI3X2),
.valid_data(TE_L1D4PHI3X1_L2D4PHI3X2_SP_L1D4PHI3X1_L2D4PHI3X2_wr_en),
.start(VMS_L2D4PHI3X2n4_start),
.done(TE_L1D4PHI3X1_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L1D4PHI3X1_L2D4PHI4X2_phi.txt","TETable_TE_L1D4PHI3X1_L2D4PHI4X2_z.txt") TE_L1D4PHI3X1_L2D4PHI4X2(
.number_in_outervmstubin(VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2_number),
.read_add_outervmstubin(VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2_read_add),
.outervmstubin(VMS_L2D4PHI4X2n2_TE_L1D4PHI3X1_L2D4PHI4X2),
.number_in_innervmstubin(VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2_number),
.read_add_innervmstubin(VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2_read_add),
.innervmstubin(VMS_L1D4PHI3X1n2_TE_L1D4PHI3X1_L2D4PHI4X2),
.stubpairout(TE_L1D4PHI3X1_L2D4PHI4X2_SP_L1D4PHI3X1_L2D4PHI4X2),
.valid_data(TE_L1D4PHI3X1_L2D4PHI4X2_SP_L1D4PHI3X1_L2D4PHI4X2_wr_en),
.start(VMS_L2D4PHI4X2n2_start),
.done(TE_L1D4PHI3X1_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI1X1_L4D3PHI1X1_phi.txt","TETable_TE_L3D3PHI1X1_L4D3PHI1X1_z.txt") TE_L3D3PHI1X1_L4D3PHI1X1(
.number_in_innervmstubin(VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_number),
.read_add_innervmstubin(VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_read_add),
.innervmstubin(VMS_L3D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1),
.number_in_outervmstubin(VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_number),
.read_add_outervmstubin(VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1_read_add),
.outervmstubin(VMS_L4D3PHI1X1n1_TE_L3D3PHI1X1_L4D3PHI1X1),
.stubpairout(TE_L3D3PHI1X1_L4D3PHI1X1_SP_L3D3PHI1X1_L4D3PHI1X1),
.valid_data(TE_L3D3PHI1X1_L4D3PHI1X1_SP_L3D3PHI1X1_L4D3PHI1X1_wr_en),
.start(VMS_L3D3PHI1X1n1_start),
.done(TE_L3D3PHI1X1_L4D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI1X1_L4D3PHI2X1_phi.txt","TETable_TE_L3D3PHI1X1_L4D3PHI2X1_z.txt") TE_L3D3PHI1X1_L4D3PHI2X1(
.number_in_innervmstubin(VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1_number),
.read_add_innervmstubin(VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1_read_add),
.innervmstubin(VMS_L3D3PHI1X1n2_TE_L3D3PHI1X1_L4D3PHI2X1),
.number_in_outervmstubin(VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1_number),
.read_add_outervmstubin(VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1_read_add),
.outervmstubin(VMS_L4D3PHI2X1n1_TE_L3D3PHI1X1_L4D3PHI2X1),
.stubpairout(TE_L3D3PHI1X1_L4D3PHI2X1_SP_L3D3PHI1X1_L4D3PHI2X1),
.valid_data(TE_L3D3PHI1X1_L4D3PHI2X1_SP_L3D3PHI1X1_L4D3PHI2X1_wr_en),
.start(VMS_L3D3PHI1X1n2_start),
.done(TE_L3D3PHI1X1_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI2X1_L4D3PHI2X1_phi.txt","TETable_TE_L3D3PHI2X1_L4D3PHI2X1_z.txt") TE_L3D3PHI2X1_L4D3PHI2X1(
.number_in_outervmstubin(VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1_number),
.read_add_outervmstubin(VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1_read_add),
.outervmstubin(VMS_L4D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI2X1),
.number_in_innervmstubin(VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1_number),
.read_add_innervmstubin(VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1_read_add),
.innervmstubin(VMS_L3D3PHI2X1n1_TE_L3D3PHI2X1_L4D3PHI2X1),
.stubpairout(TE_L3D3PHI2X1_L4D3PHI2X1_SP_L3D3PHI2X1_L4D3PHI2X1),
.valid_data(TE_L3D3PHI2X1_L4D3PHI2X1_SP_L3D3PHI2X1_L4D3PHI2X1_wr_en),
.start(VMS_L4D3PHI2X1n2_start),
.done(TE_L3D3PHI2X1_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI2X1_L4D3PHI3X1_phi.txt","TETable_TE_L3D3PHI2X1_L4D3PHI3X1_z.txt") TE_L3D3PHI2X1_L4D3PHI3X1(
.number_in_innervmstubin(VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1_number),
.read_add_innervmstubin(VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1_read_add),
.innervmstubin(VMS_L3D3PHI2X1n2_TE_L3D3PHI2X1_L4D3PHI3X1),
.number_in_outervmstubin(VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1_number),
.read_add_outervmstubin(VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1_read_add),
.outervmstubin(VMS_L4D3PHI3X1n1_TE_L3D3PHI2X1_L4D3PHI3X1),
.stubpairout(TE_L3D3PHI2X1_L4D3PHI3X1_SP_L3D3PHI2X1_L4D3PHI3X1),
.valid_data(TE_L3D3PHI2X1_L4D3PHI3X1_SP_L3D3PHI2X1_L4D3PHI3X1_wr_en),
.start(VMS_L3D3PHI2X1n2_start),
.done(TE_L3D3PHI2X1_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI3X1_L4D3PHI3X1_phi.txt","TETable_TE_L3D3PHI3X1_L4D3PHI3X1_z.txt") TE_L3D3PHI3X1_L4D3PHI3X1(
.number_in_outervmstubin(VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1_number),
.read_add_outervmstubin(VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1_read_add),
.outervmstubin(VMS_L4D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI3X1),
.number_in_innervmstubin(VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1_number),
.read_add_innervmstubin(VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1_read_add),
.innervmstubin(VMS_L3D3PHI3X1n1_TE_L3D3PHI3X1_L4D3PHI3X1),
.stubpairout(TE_L3D3PHI3X1_L4D3PHI3X1_SP_L3D3PHI3X1_L4D3PHI3X1),
.valid_data(TE_L3D3PHI3X1_L4D3PHI3X1_SP_L3D3PHI3X1_L4D3PHI3X1_wr_en),
.start(VMS_L4D3PHI3X1n2_start),
.done(TE_L3D3PHI3X1_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI3X1_L4D3PHI4X1_phi.txt","TETable_TE_L3D3PHI3X1_L4D3PHI4X1_z.txt") TE_L3D3PHI3X1_L4D3PHI4X1(
.number_in_innervmstubin(VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1_number),
.read_add_innervmstubin(VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1_read_add),
.innervmstubin(VMS_L3D3PHI3X1n2_TE_L3D3PHI3X1_L4D3PHI4X1),
.number_in_outervmstubin(VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1_number),
.read_add_outervmstubin(VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1_read_add),
.outervmstubin(VMS_L4D3PHI4X1n1_TE_L3D3PHI3X1_L4D3PHI4X1),
.stubpairout(TE_L3D3PHI3X1_L4D3PHI4X1_SP_L3D3PHI3X1_L4D3PHI4X1),
.valid_data(TE_L3D3PHI3X1_L4D3PHI4X1_SP_L3D3PHI3X1_L4D3PHI4X1_wr_en),
.start(VMS_L3D3PHI3X1n2_start),
.done(TE_L3D3PHI3X1_L4D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI1X2_L4D3PHI1X2_phi.txt","TETable_TE_L3D3PHI1X2_L4D3PHI1X2_z.txt") TE_L3D3PHI1X2_L4D3PHI1X2(
.number_in_innervmstubin(VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_number),
.read_add_innervmstubin(VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_read_add),
.innervmstubin(VMS_L3D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2),
.number_in_outervmstubin(VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_number),
.read_add_outervmstubin(VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2_read_add),
.outervmstubin(VMS_L4D3PHI1X2n1_TE_L3D3PHI1X2_L4D3PHI1X2),
.stubpairout(TE_L3D3PHI1X2_L4D3PHI1X2_SP_L3D3PHI1X2_L4D3PHI1X2),
.valid_data(TE_L3D3PHI1X2_L4D3PHI1X2_SP_L3D3PHI1X2_L4D3PHI1X2_wr_en),
.start(VMS_L3D3PHI1X2n1_start),
.done(TE_L3D3PHI1X2_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI1X2_L4D3PHI2X2_phi.txt","TETable_TE_L3D3PHI1X2_L4D3PHI2X2_z.txt") TE_L3D3PHI1X2_L4D3PHI2X2(
.number_in_innervmstubin(VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2_number),
.read_add_innervmstubin(VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2_read_add),
.innervmstubin(VMS_L3D3PHI1X2n2_TE_L3D3PHI1X2_L4D3PHI2X2),
.number_in_outervmstubin(VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2_number),
.read_add_outervmstubin(VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2_read_add),
.outervmstubin(VMS_L4D3PHI2X2n1_TE_L3D3PHI1X2_L4D3PHI2X2),
.stubpairout(TE_L3D3PHI1X2_L4D3PHI2X2_SP_L3D3PHI1X2_L4D3PHI2X2),
.valid_data(TE_L3D3PHI1X2_L4D3PHI2X2_SP_L3D3PHI1X2_L4D3PHI2X2_wr_en),
.start(VMS_L3D3PHI1X2n2_start),
.done(TE_L3D3PHI1X2_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI2X2_L4D3PHI2X2_phi.txt","TETable_TE_L3D3PHI2X2_L4D3PHI2X2_z.txt") TE_L3D3PHI2X2_L4D3PHI2X2(
.number_in_outervmstubin(VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2_number),
.read_add_outervmstubin(VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2_read_add),
.outervmstubin(VMS_L4D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI2X2),
.number_in_innervmstubin(VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2_number),
.read_add_innervmstubin(VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2_read_add),
.innervmstubin(VMS_L3D3PHI2X2n1_TE_L3D3PHI2X2_L4D3PHI2X2),
.stubpairout(TE_L3D3PHI2X2_L4D3PHI2X2_SP_L3D3PHI2X2_L4D3PHI2X2),
.valid_data(TE_L3D3PHI2X2_L4D3PHI2X2_SP_L3D3PHI2X2_L4D3PHI2X2_wr_en),
.start(VMS_L4D3PHI2X2n2_start),
.done(TE_L3D3PHI2X2_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI2X2_L4D3PHI3X2_phi.txt","TETable_TE_L3D3PHI2X2_L4D3PHI3X2_z.txt") TE_L3D3PHI2X2_L4D3PHI3X2(
.number_in_innervmstubin(VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2_number),
.read_add_innervmstubin(VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2_read_add),
.innervmstubin(VMS_L3D3PHI2X2n2_TE_L3D3PHI2X2_L4D3PHI3X2),
.number_in_outervmstubin(VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2_number),
.read_add_outervmstubin(VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2_read_add),
.outervmstubin(VMS_L4D3PHI3X2n1_TE_L3D3PHI2X2_L4D3PHI3X2),
.stubpairout(TE_L3D3PHI2X2_L4D3PHI3X2_SP_L3D3PHI2X2_L4D3PHI3X2),
.valid_data(TE_L3D3PHI2X2_L4D3PHI3X2_SP_L3D3PHI2X2_L4D3PHI3X2_wr_en),
.start(VMS_L3D3PHI2X2n2_start),
.done(TE_L3D3PHI2X2_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI3X2_L4D3PHI3X2_phi.txt","TETable_TE_L3D3PHI3X2_L4D3PHI3X2_z.txt") TE_L3D3PHI3X2_L4D3PHI3X2(
.number_in_outervmstubin(VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2_number),
.read_add_outervmstubin(VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2_read_add),
.outervmstubin(VMS_L4D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI3X2),
.number_in_innervmstubin(VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2_number),
.read_add_innervmstubin(VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2_read_add),
.innervmstubin(VMS_L3D3PHI3X2n1_TE_L3D3PHI3X2_L4D3PHI3X2),
.stubpairout(TE_L3D3PHI3X2_L4D3PHI3X2_SP_L3D3PHI3X2_L4D3PHI3X2),
.valid_data(TE_L3D3PHI3X2_L4D3PHI3X2_SP_L3D3PHI3X2_L4D3PHI3X2_wr_en),
.start(VMS_L4D3PHI3X2n2_start),
.done(TE_L3D3PHI3X2_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI3X2_L4D3PHI4X2_phi.txt","TETable_TE_L3D3PHI3X2_L4D3PHI4X2_z.txt") TE_L3D3PHI3X2_L4D3PHI4X2(
.number_in_innervmstubin(VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2_number),
.read_add_innervmstubin(VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2_read_add),
.innervmstubin(VMS_L3D3PHI3X2n2_TE_L3D3PHI3X2_L4D3PHI4X2),
.number_in_outervmstubin(VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2_number),
.read_add_outervmstubin(VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2_read_add),
.outervmstubin(VMS_L4D3PHI4X2n1_TE_L3D3PHI3X2_L4D3PHI4X2),
.stubpairout(TE_L3D3PHI3X2_L4D3PHI4X2_SP_L3D3PHI3X2_L4D3PHI4X2),
.valid_data(TE_L3D3PHI3X2_L4D3PHI4X2_SP_L3D3PHI3X2_L4D3PHI4X2_wr_en),
.start(VMS_L3D3PHI3X2n2_start),
.done(TE_L3D3PHI3X2_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI1X1_L4D3PHI1X2_phi.txt","TETable_TE_L3D3PHI1X1_L4D3PHI1X2_z.txt") TE_L3D3PHI1X1_L4D3PHI1X2(
.number_in_innervmstubin(VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2_number),
.read_add_innervmstubin(VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2_read_add),
.innervmstubin(VMS_L3D3PHI1X1n3_TE_L3D3PHI1X1_L4D3PHI1X2),
.number_in_outervmstubin(VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2_number),
.read_add_outervmstubin(VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2_read_add),
.outervmstubin(VMS_L4D3PHI1X2n2_TE_L3D3PHI1X1_L4D3PHI1X2),
.stubpairout(TE_L3D3PHI1X1_L4D3PHI1X2_SP_L3D3PHI1X1_L4D3PHI1X2),
.valid_data(TE_L3D3PHI1X1_L4D3PHI1X2_SP_L3D3PHI1X1_L4D3PHI1X2_wr_en),
.start(VMS_L3D3PHI1X1n3_start),
.done(TE_L3D3PHI1X1_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI1X1_L4D3PHI2X2_phi.txt","TETable_TE_L3D3PHI1X1_L4D3PHI2X2_z.txt") TE_L3D3PHI1X1_L4D3PHI2X2(
.number_in_innervmstubin(VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2_number),
.read_add_innervmstubin(VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2_read_add),
.innervmstubin(VMS_L3D3PHI1X1n4_TE_L3D3PHI1X1_L4D3PHI2X2),
.number_in_outervmstubin(VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2_number),
.read_add_outervmstubin(VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2_read_add),
.outervmstubin(VMS_L4D3PHI2X2n3_TE_L3D3PHI1X1_L4D3PHI2X2),
.stubpairout(TE_L3D3PHI1X1_L4D3PHI2X2_SP_L3D3PHI1X1_L4D3PHI2X2),
.valid_data(TE_L3D3PHI1X1_L4D3PHI2X2_SP_L3D3PHI1X1_L4D3PHI2X2_wr_en),
.start(VMS_L3D3PHI1X1n4_start),
.done(TE_L3D3PHI1X1_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI2X1_L4D3PHI2X2_phi.txt","TETable_TE_L3D3PHI2X1_L4D3PHI2X2_z.txt") TE_L3D3PHI2X1_L4D3PHI2X2(
.number_in_innervmstubin(VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2_number),
.read_add_innervmstubin(VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2_read_add),
.innervmstubin(VMS_L3D3PHI2X1n3_TE_L3D3PHI2X1_L4D3PHI2X2),
.number_in_outervmstubin(VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2_number),
.read_add_outervmstubin(VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2_read_add),
.outervmstubin(VMS_L4D3PHI2X2n4_TE_L3D3PHI2X1_L4D3PHI2X2),
.stubpairout(TE_L3D3PHI2X1_L4D3PHI2X2_SP_L3D3PHI2X1_L4D3PHI2X2),
.valid_data(TE_L3D3PHI2X1_L4D3PHI2X2_SP_L3D3PHI2X1_L4D3PHI2X2_wr_en),
.start(VMS_L3D3PHI2X1n3_start),
.done(TE_L3D3PHI2X1_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI2X1_L4D3PHI3X2_phi.txt","TETable_TE_L3D3PHI2X1_L4D3PHI3X2_z.txt") TE_L3D3PHI2X1_L4D3PHI3X2(
.number_in_innervmstubin(VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2_number),
.read_add_innervmstubin(VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2_read_add),
.innervmstubin(VMS_L3D3PHI2X1n4_TE_L3D3PHI2X1_L4D3PHI3X2),
.number_in_outervmstubin(VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2_number),
.read_add_outervmstubin(VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2_read_add),
.outervmstubin(VMS_L4D3PHI3X2n3_TE_L3D3PHI2X1_L4D3PHI3X2),
.stubpairout(TE_L3D3PHI2X1_L4D3PHI3X2_SP_L3D3PHI2X1_L4D3PHI3X2),
.valid_data(TE_L3D3PHI2X1_L4D3PHI3X2_SP_L3D3PHI2X1_L4D3PHI3X2_wr_en),
.start(VMS_L3D3PHI2X1n4_start),
.done(TE_L3D3PHI2X1_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI3X1_L4D3PHI3X2_phi.txt","TETable_TE_L3D3PHI3X1_L4D3PHI3X2_z.txt") TE_L3D3PHI3X1_L4D3PHI3X2(
.number_in_innervmstubin(VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2_number),
.read_add_innervmstubin(VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2_read_add),
.innervmstubin(VMS_L3D3PHI3X1n3_TE_L3D3PHI3X1_L4D3PHI3X2),
.number_in_outervmstubin(VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2_number),
.read_add_outervmstubin(VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2_read_add),
.outervmstubin(VMS_L4D3PHI3X2n4_TE_L3D3PHI3X1_L4D3PHI3X2),
.stubpairout(TE_L3D3PHI3X1_L4D3PHI3X2_SP_L3D3PHI3X1_L4D3PHI3X2),
.valid_data(TE_L3D3PHI3X1_L4D3PHI3X2_SP_L3D3PHI3X1_L4D3PHI3X2_wr_en),
.start(VMS_L3D3PHI3X1n3_start),
.done(TE_L3D3PHI3X1_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI3X1_L4D3PHI4X2_phi.txt","TETable_TE_L3D3PHI3X1_L4D3PHI4X2_z.txt") TE_L3D3PHI3X1_L4D3PHI4X2(
.number_in_innervmstubin(VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2_number),
.read_add_innervmstubin(VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2_read_add),
.innervmstubin(VMS_L3D3PHI3X1n4_TE_L3D3PHI3X1_L4D3PHI4X2),
.number_in_outervmstubin(VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2_number),
.read_add_outervmstubin(VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2_read_add),
.outervmstubin(VMS_L4D3PHI4X2n2_TE_L3D3PHI3X1_L4D3PHI4X2),
.stubpairout(TE_L3D3PHI3X1_L4D3PHI4X2_SP_L3D3PHI3X1_L4D3PHI4X2),
.valid_data(TE_L3D3PHI3X1_L4D3PHI4X2_SP_L3D3PHI3X1_L4D3PHI4X2_wr_en),
.start(VMS_L3D3PHI3X1n4_start),
.done(TE_L3D3PHI3X1_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI1X2_L4D4PHI1X1_phi.txt","TETable_TE_L3D3PHI1X2_L4D4PHI1X1_z.txt") TE_L3D3PHI1X2_L4D4PHI1X1(
.number_in_innervmstubin(VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1_number),
.read_add_innervmstubin(VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1_read_add),
.innervmstubin(VMS_L3D3PHI1X2n3_TE_L3D3PHI1X2_L4D4PHI1X1),
.number_in_outervmstubin(VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1_number),
.read_add_outervmstubin(VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1_read_add),
.outervmstubin(VMS_L4D4PHI1X1n1_TE_L3D3PHI1X2_L4D4PHI1X1),
.stubpairout(TE_L3D3PHI1X2_L4D4PHI1X1_SP_L3D3PHI1X2_L4D4PHI1X1),
.valid_data(TE_L3D3PHI1X2_L4D4PHI1X1_SP_L3D3PHI1X2_L4D4PHI1X1_wr_en),
.start(VMS_L3D3PHI1X2n3_start),
.done(TE_L3D3PHI1X2_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI1X2_L4D4PHI2X1_phi.txt","TETable_TE_L3D3PHI1X2_L4D4PHI2X1_z.txt") TE_L3D3PHI1X2_L4D4PHI2X1(
.number_in_innervmstubin(VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1_number),
.read_add_innervmstubin(VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1_read_add),
.innervmstubin(VMS_L3D3PHI1X2n4_TE_L3D3PHI1X2_L4D4PHI2X1),
.number_in_outervmstubin(VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1_number),
.read_add_outervmstubin(VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1_read_add),
.outervmstubin(VMS_L4D4PHI2X1n1_TE_L3D3PHI1X2_L4D4PHI2X1),
.stubpairout(TE_L3D3PHI1X2_L4D4PHI2X1_SP_L3D3PHI1X2_L4D4PHI2X1),
.valid_data(TE_L3D3PHI1X2_L4D4PHI2X1_SP_L3D3PHI1X2_L4D4PHI2X1_wr_en),
.start(VMS_L3D3PHI1X2n4_start),
.done(TE_L3D3PHI1X2_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI2X2_L4D4PHI2X1_phi.txt","TETable_TE_L3D3PHI2X2_L4D4PHI2X1_z.txt") TE_L3D3PHI2X2_L4D4PHI2X1(
.number_in_innervmstubin(VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1_number),
.read_add_innervmstubin(VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1_read_add),
.innervmstubin(VMS_L3D3PHI2X2n3_TE_L3D3PHI2X2_L4D4PHI2X1),
.number_in_outervmstubin(VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1_number),
.read_add_outervmstubin(VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1_read_add),
.outervmstubin(VMS_L4D4PHI2X1n2_TE_L3D3PHI2X2_L4D4PHI2X1),
.stubpairout(TE_L3D3PHI2X2_L4D4PHI2X1_SP_L3D3PHI2X2_L4D4PHI2X1),
.valid_data(TE_L3D3PHI2X2_L4D4PHI2X1_SP_L3D3PHI2X2_L4D4PHI2X1_wr_en),
.start(VMS_L3D3PHI2X2n3_start),
.done(TE_L3D3PHI2X2_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI2X2_L4D4PHI3X1_phi.txt","TETable_TE_L3D3PHI2X2_L4D4PHI3X1_z.txt") TE_L3D3PHI2X2_L4D4PHI3X1(
.number_in_innervmstubin(VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1_number),
.read_add_innervmstubin(VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1_read_add),
.innervmstubin(VMS_L3D3PHI2X2n4_TE_L3D3PHI2X2_L4D4PHI3X1),
.number_in_outervmstubin(VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1_number),
.read_add_outervmstubin(VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1_read_add),
.outervmstubin(VMS_L4D4PHI3X1n1_TE_L3D3PHI2X2_L4D4PHI3X1),
.stubpairout(TE_L3D3PHI2X2_L4D4PHI3X1_SP_L3D3PHI2X2_L4D4PHI3X1),
.valid_data(TE_L3D3PHI2X2_L4D4PHI3X1_SP_L3D3PHI2X2_L4D4PHI3X1_wr_en),
.start(VMS_L3D3PHI2X2n4_start),
.done(TE_L3D3PHI2X2_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI3X2_L4D4PHI3X1_phi.txt","TETable_TE_L3D3PHI3X2_L4D4PHI3X1_z.txt") TE_L3D3PHI3X2_L4D4PHI3X1(
.number_in_innervmstubin(VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1_number),
.read_add_innervmstubin(VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1_read_add),
.innervmstubin(VMS_L3D3PHI3X2n3_TE_L3D3PHI3X2_L4D4PHI3X1),
.number_in_outervmstubin(VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1_number),
.read_add_outervmstubin(VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1_read_add),
.outervmstubin(VMS_L4D4PHI3X1n2_TE_L3D3PHI3X2_L4D4PHI3X1),
.stubpairout(TE_L3D3PHI3X2_L4D4PHI3X1_SP_L3D3PHI3X2_L4D4PHI3X1),
.valid_data(TE_L3D3PHI3X2_L4D4PHI3X1_SP_L3D3PHI3X2_L4D4PHI3X1_wr_en),
.start(VMS_L3D3PHI3X2n3_start),
.done(TE_L3D3PHI3X2_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D3PHI3X2_L4D4PHI4X1_phi.txt","TETable_TE_L3D3PHI3X2_L4D4PHI4X1_z.txt") TE_L3D3PHI3X2_L4D4PHI4X1(
.number_in_innervmstubin(VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1_number),
.read_add_innervmstubin(VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1_read_add),
.innervmstubin(VMS_L3D3PHI3X2n4_TE_L3D3PHI3X2_L4D4PHI4X1),
.number_in_outervmstubin(VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1_number),
.read_add_outervmstubin(VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1_read_add),
.outervmstubin(VMS_L4D4PHI4X1n1_TE_L3D3PHI3X2_L4D4PHI4X1),
.stubpairout(TE_L3D3PHI3X2_L4D4PHI4X1_SP_L3D3PHI3X2_L4D4PHI4X1),
.valid_data(TE_L3D3PHI3X2_L4D4PHI4X1_SP_L3D3PHI3X2_L4D4PHI4X1_wr_en),
.start(VMS_L3D3PHI3X2n4_start),
.done(TE_L3D3PHI3X2_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI1X1_L4D4PHI1X1_phi.txt","TETable_TE_L3D4PHI1X1_L4D4PHI1X1_z.txt") TE_L3D4PHI1X1_L4D4PHI1X1(
.number_in_outervmstubin(VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1_number),
.read_add_outervmstubin(VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1_read_add),
.outervmstubin(VMS_L4D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI1X1),
.number_in_innervmstubin(VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1_number),
.read_add_innervmstubin(VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1_read_add),
.innervmstubin(VMS_L3D4PHI1X1n1_TE_L3D4PHI1X1_L4D4PHI1X1),
.stubpairout(TE_L3D4PHI1X1_L4D4PHI1X1_SP_L3D4PHI1X1_L4D4PHI1X1),
.valid_data(TE_L3D4PHI1X1_L4D4PHI1X1_SP_L3D4PHI1X1_L4D4PHI1X1_wr_en),
.start(VMS_L4D4PHI1X1n2_start),
.done(TE_L3D4PHI1X1_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI1X1_L4D4PHI2X1_phi.txt","TETable_TE_L3D4PHI1X1_L4D4PHI2X1_z.txt") TE_L3D4PHI1X1_L4D4PHI2X1(
.number_in_outervmstubin(VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1_number),
.read_add_outervmstubin(VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1_read_add),
.outervmstubin(VMS_L4D4PHI2X1n3_TE_L3D4PHI1X1_L4D4PHI2X1),
.number_in_innervmstubin(VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1_number),
.read_add_innervmstubin(VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1_read_add),
.innervmstubin(VMS_L3D4PHI1X1n2_TE_L3D4PHI1X1_L4D4PHI2X1),
.stubpairout(TE_L3D4PHI1X1_L4D4PHI2X1_SP_L3D4PHI1X1_L4D4PHI2X1),
.valid_data(TE_L3D4PHI1X1_L4D4PHI2X1_SP_L3D4PHI1X1_L4D4PHI2X1_wr_en),
.start(VMS_L4D4PHI2X1n3_start),
.done(TE_L3D4PHI1X1_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI2X1_L4D4PHI2X1_phi.txt","TETable_TE_L3D4PHI2X1_L4D4PHI2X1_z.txt") TE_L3D4PHI2X1_L4D4PHI2X1(
.number_in_outervmstubin(VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1_number),
.read_add_outervmstubin(VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1_read_add),
.outervmstubin(VMS_L4D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI2X1),
.number_in_innervmstubin(VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1_number),
.read_add_innervmstubin(VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1_read_add),
.innervmstubin(VMS_L3D4PHI2X1n1_TE_L3D4PHI2X1_L4D4PHI2X1),
.stubpairout(TE_L3D4PHI2X1_L4D4PHI2X1_SP_L3D4PHI2X1_L4D4PHI2X1),
.valid_data(TE_L3D4PHI2X1_L4D4PHI2X1_SP_L3D4PHI2X1_L4D4PHI2X1_wr_en),
.start(VMS_L4D4PHI2X1n4_start),
.done(TE_L3D4PHI2X1_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI2X1_L4D4PHI3X1_phi.txt","TETable_TE_L3D4PHI2X1_L4D4PHI3X1_z.txt") TE_L3D4PHI2X1_L4D4PHI3X1(
.number_in_outervmstubin(VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1_number),
.read_add_outervmstubin(VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1_read_add),
.outervmstubin(VMS_L4D4PHI3X1n3_TE_L3D4PHI2X1_L4D4PHI3X1),
.number_in_innervmstubin(VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1_number),
.read_add_innervmstubin(VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1_read_add),
.innervmstubin(VMS_L3D4PHI2X1n2_TE_L3D4PHI2X1_L4D4PHI3X1),
.stubpairout(TE_L3D4PHI2X1_L4D4PHI3X1_SP_L3D4PHI2X1_L4D4PHI3X1),
.valid_data(TE_L3D4PHI2X1_L4D4PHI3X1_SP_L3D4PHI2X1_L4D4PHI3X1_wr_en),
.start(VMS_L4D4PHI3X1n3_start),
.done(TE_L3D4PHI2X1_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI3X1_L4D4PHI3X1_phi.txt","TETable_TE_L3D4PHI3X1_L4D4PHI3X1_z.txt") TE_L3D4PHI3X1_L4D4PHI3X1(
.number_in_outervmstubin(VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1_number),
.read_add_outervmstubin(VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1_read_add),
.outervmstubin(VMS_L4D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI3X1),
.number_in_innervmstubin(VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1_number),
.read_add_innervmstubin(VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1_read_add),
.innervmstubin(VMS_L3D4PHI3X1n1_TE_L3D4PHI3X1_L4D4PHI3X1),
.stubpairout(TE_L3D4PHI3X1_L4D4PHI3X1_SP_L3D4PHI3X1_L4D4PHI3X1),
.valid_data(TE_L3D4PHI3X1_L4D4PHI3X1_SP_L3D4PHI3X1_L4D4PHI3X1_wr_en),
.start(VMS_L4D4PHI3X1n4_start),
.done(TE_L3D4PHI3X1_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI3X1_L4D4PHI4X1_phi.txt","TETable_TE_L3D4PHI3X1_L4D4PHI4X1_z.txt") TE_L3D4PHI3X1_L4D4PHI4X1(
.number_in_outervmstubin(VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_number),
.read_add_outervmstubin(VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_read_add),
.outervmstubin(VMS_L4D4PHI4X1n2_TE_L3D4PHI3X1_L4D4PHI4X1),
.number_in_innervmstubin(VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_number),
.read_add_innervmstubin(VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1_read_add),
.innervmstubin(VMS_L3D4PHI3X1n2_TE_L3D4PHI3X1_L4D4PHI4X1),
.stubpairout(TE_L3D4PHI3X1_L4D4PHI4X1_SP_L3D4PHI3X1_L4D4PHI4X1),
.valid_data(TE_L3D4PHI3X1_L4D4PHI4X1_SP_L3D4PHI3X1_L4D4PHI4X1_wr_en),
.start(VMS_L4D4PHI4X1n2_start),
.done(TE_L3D4PHI3X1_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI1X1_L4D4PHI1X2_phi.txt","TETable_TE_L3D4PHI1X1_L4D4PHI1X2_z.txt") TE_L3D4PHI1X1_L4D4PHI1X2(
.number_in_innervmstubin(VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2_number),
.read_add_innervmstubin(VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2_read_add),
.innervmstubin(VMS_L3D4PHI1X1n3_TE_L3D4PHI1X1_L4D4PHI1X2),
.number_in_outervmstubin(VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2_number),
.read_add_outervmstubin(VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2_read_add),
.outervmstubin(VMS_L4D4PHI1X2n1_TE_L3D4PHI1X1_L4D4PHI1X2),
.stubpairout(TE_L3D4PHI1X1_L4D4PHI1X2_SP_L3D4PHI1X1_L4D4PHI1X2),
.valid_data(TE_L3D4PHI1X1_L4D4PHI1X2_SP_L3D4PHI1X1_L4D4PHI1X2_wr_en),
.start(VMS_L3D4PHI1X1n3_start),
.done(TE_L3D4PHI1X1_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI1X1_L4D4PHI2X2_phi.txt","TETable_TE_L3D4PHI1X1_L4D4PHI2X2_z.txt") TE_L3D4PHI1X1_L4D4PHI2X2(
.number_in_innervmstubin(VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2_number),
.read_add_innervmstubin(VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2_read_add),
.innervmstubin(VMS_L3D4PHI1X1n4_TE_L3D4PHI1X1_L4D4PHI2X2),
.number_in_outervmstubin(VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2_number),
.read_add_outervmstubin(VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2_read_add),
.outervmstubin(VMS_L4D4PHI2X2n1_TE_L3D4PHI1X1_L4D4PHI2X2),
.stubpairout(TE_L3D4PHI1X1_L4D4PHI2X2_SP_L3D4PHI1X1_L4D4PHI2X2),
.valid_data(TE_L3D4PHI1X1_L4D4PHI2X2_SP_L3D4PHI1X1_L4D4PHI2X2_wr_en),
.start(VMS_L3D4PHI1X1n4_start),
.done(TE_L3D4PHI1X1_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI2X1_L4D4PHI2X2_phi.txt","TETable_TE_L3D4PHI2X1_L4D4PHI2X2_z.txt") TE_L3D4PHI2X1_L4D4PHI2X2(
.number_in_innervmstubin(VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2_number),
.read_add_innervmstubin(VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2_read_add),
.innervmstubin(VMS_L3D4PHI2X1n3_TE_L3D4PHI2X1_L4D4PHI2X2),
.number_in_outervmstubin(VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2_number),
.read_add_outervmstubin(VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2_read_add),
.outervmstubin(VMS_L4D4PHI2X2n2_TE_L3D4PHI2X1_L4D4PHI2X2),
.stubpairout(TE_L3D4PHI2X1_L4D4PHI2X2_SP_L3D4PHI2X1_L4D4PHI2X2),
.valid_data(TE_L3D4PHI2X1_L4D4PHI2X2_SP_L3D4PHI2X1_L4D4PHI2X2_wr_en),
.start(VMS_L3D4PHI2X1n3_start),
.done(TE_L3D4PHI2X1_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI2X1_L4D4PHI3X2_phi.txt","TETable_TE_L3D4PHI2X1_L4D4PHI3X2_z.txt") TE_L3D4PHI2X1_L4D4PHI3X2(
.number_in_innervmstubin(VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2_number),
.read_add_innervmstubin(VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2_read_add),
.innervmstubin(VMS_L3D4PHI2X1n4_TE_L3D4PHI2X1_L4D4PHI3X2),
.number_in_outervmstubin(VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2_number),
.read_add_outervmstubin(VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2_read_add),
.outervmstubin(VMS_L4D4PHI3X2n1_TE_L3D4PHI2X1_L4D4PHI3X2),
.stubpairout(TE_L3D4PHI2X1_L4D4PHI3X2_SP_L3D4PHI2X1_L4D4PHI3X2),
.valid_data(TE_L3D4PHI2X1_L4D4PHI3X2_SP_L3D4PHI2X1_L4D4PHI3X2_wr_en),
.start(VMS_L3D4PHI2X1n4_start),
.done(TE_L3D4PHI2X1_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI3X1_L4D4PHI3X2_phi.txt","TETable_TE_L3D4PHI3X1_L4D4PHI3X2_z.txt") TE_L3D4PHI3X1_L4D4PHI3X2(
.number_in_innervmstubin(VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2_number),
.read_add_innervmstubin(VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2_read_add),
.innervmstubin(VMS_L3D4PHI3X1n3_TE_L3D4PHI3X1_L4D4PHI3X2),
.number_in_outervmstubin(VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2_number),
.read_add_outervmstubin(VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2_read_add),
.outervmstubin(VMS_L4D4PHI3X2n2_TE_L3D4PHI3X1_L4D4PHI3X2),
.stubpairout(TE_L3D4PHI3X1_L4D4PHI3X2_SP_L3D4PHI3X1_L4D4PHI3X2),
.valid_data(TE_L3D4PHI3X1_L4D4PHI3X2_SP_L3D4PHI3X1_L4D4PHI3X2_wr_en),
.start(VMS_L3D4PHI3X1n3_start),
.done(TE_L3D4PHI3X1_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI3X1_L4D4PHI4X2_phi.txt","TETable_TE_L3D4PHI3X1_L4D4PHI4X2_z.txt") TE_L3D4PHI3X1_L4D4PHI4X2(
.number_in_innervmstubin(VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2_number),
.read_add_innervmstubin(VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2_read_add),
.innervmstubin(VMS_L3D4PHI3X1n4_TE_L3D4PHI3X1_L4D4PHI4X2),
.number_in_outervmstubin(VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2_number),
.read_add_outervmstubin(VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2_read_add),
.outervmstubin(VMS_L4D4PHI4X2n1_TE_L3D4PHI3X1_L4D4PHI4X2),
.stubpairout(TE_L3D4PHI3X1_L4D4PHI4X2_SP_L3D4PHI3X1_L4D4PHI4X2),
.valid_data(TE_L3D4PHI3X1_L4D4PHI4X2_SP_L3D4PHI3X1_L4D4PHI4X2_wr_en),
.start(VMS_L3D4PHI3X1n4_start),
.done(TE_L3D4PHI3X1_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI1X2_L4D4PHI1X2_phi.txt","TETable_TE_L3D4PHI1X2_L4D4PHI1X2_z.txt") TE_L3D4PHI1X2_L4D4PHI1X2(
.number_in_outervmstubin(VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2_number),
.read_add_outervmstubin(VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2_read_add),
.outervmstubin(VMS_L4D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI1X2),
.number_in_innervmstubin(VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2_number),
.read_add_innervmstubin(VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2_read_add),
.innervmstubin(VMS_L3D4PHI1X2n1_TE_L3D4PHI1X2_L4D4PHI1X2),
.stubpairout(TE_L3D4PHI1X2_L4D4PHI1X2_SP_L3D4PHI1X2_L4D4PHI1X2),
.valid_data(TE_L3D4PHI1X2_L4D4PHI1X2_SP_L3D4PHI1X2_L4D4PHI1X2_wr_en),
.start(VMS_L4D4PHI1X2n2_start),
.done(TE_L3D4PHI1X2_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI1X2_L4D4PHI2X2_phi.txt","TETable_TE_L3D4PHI1X2_L4D4PHI2X2_z.txt") TE_L3D4PHI1X2_L4D4PHI2X2(
.number_in_outervmstubin(VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2_number),
.read_add_outervmstubin(VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2_read_add),
.outervmstubin(VMS_L4D4PHI2X2n3_TE_L3D4PHI1X2_L4D4PHI2X2),
.number_in_innervmstubin(VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2_number),
.read_add_innervmstubin(VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2_read_add),
.innervmstubin(VMS_L3D4PHI1X2n2_TE_L3D4PHI1X2_L4D4PHI2X2),
.stubpairout(TE_L3D4PHI1X2_L4D4PHI2X2_SP_L3D4PHI1X2_L4D4PHI2X2),
.valid_data(TE_L3D4PHI1X2_L4D4PHI2X2_SP_L3D4PHI1X2_L4D4PHI2X2_wr_en),
.start(VMS_L4D4PHI2X2n3_start),
.done(TE_L3D4PHI1X2_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI2X2_L4D4PHI2X2_phi.txt","TETable_TE_L3D4PHI2X2_L4D4PHI2X2_z.txt") TE_L3D4PHI2X2_L4D4PHI2X2(
.number_in_outervmstubin(VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2_number),
.read_add_outervmstubin(VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2_read_add),
.outervmstubin(VMS_L4D4PHI2X2n4_TE_L3D4PHI2X2_L4D4PHI2X2),
.number_in_innervmstubin(VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2_number),
.read_add_innervmstubin(VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2_read_add),
.innervmstubin(VMS_L3D4PHI2X2n1_TE_L3D4PHI2X2_L4D4PHI2X2),
.stubpairout(TE_L3D4PHI2X2_L4D4PHI2X2_SP_L3D4PHI2X2_L4D4PHI2X2),
.valid_data(TE_L3D4PHI2X2_L4D4PHI2X2_SP_L3D4PHI2X2_L4D4PHI2X2_wr_en),
.start(VMS_L4D4PHI2X2n4_start),
.done(TE_L3D4PHI2X2_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI2X2_L4D4PHI3X2_phi.txt","TETable_TE_L3D4PHI2X2_L4D4PHI3X2_z.txt") TE_L3D4PHI2X2_L4D4PHI3X2(
.number_in_outervmstubin(VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2_number),
.read_add_outervmstubin(VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2_read_add),
.outervmstubin(VMS_L4D4PHI3X2n3_TE_L3D4PHI2X2_L4D4PHI3X2),
.number_in_innervmstubin(VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2_number),
.read_add_innervmstubin(VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2_read_add),
.innervmstubin(VMS_L3D4PHI2X2n2_TE_L3D4PHI2X2_L4D4PHI3X2),
.stubpairout(TE_L3D4PHI2X2_L4D4PHI3X2_SP_L3D4PHI2X2_L4D4PHI3X2),
.valid_data(TE_L3D4PHI2X2_L4D4PHI3X2_SP_L3D4PHI2X2_L4D4PHI3X2_wr_en),
.start(VMS_L4D4PHI3X2n3_start),
.done(TE_L3D4PHI2X2_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI3X2_L4D4PHI3X2_phi.txt","TETable_TE_L3D4PHI3X2_L4D4PHI3X2_z.txt") TE_L3D4PHI3X2_L4D4PHI3X2(
.number_in_outervmstubin(VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2_number),
.read_add_outervmstubin(VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2_read_add),
.outervmstubin(VMS_L4D4PHI3X2n4_TE_L3D4PHI3X2_L4D4PHI3X2),
.number_in_innervmstubin(VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2_number),
.read_add_innervmstubin(VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2_read_add),
.innervmstubin(VMS_L3D4PHI3X2n1_TE_L3D4PHI3X2_L4D4PHI3X2),
.stubpairout(TE_L3D4PHI3X2_L4D4PHI3X2_SP_L3D4PHI3X2_L4D4PHI3X2),
.valid_data(TE_L3D4PHI3X2_L4D4PHI3X2_SP_L3D4PHI3X2_L4D4PHI3X2_wr_en),
.start(VMS_L4D4PHI3X2n4_start),
.done(TE_L3D4PHI3X2_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L3D4PHI3X2_L4D4PHI4X2_phi.txt","TETable_TE_L3D4PHI3X2_L4D4PHI4X2_z.txt") TE_L3D4PHI3X2_L4D4PHI4X2(
.number_in_outervmstubin(VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_number),
.read_add_outervmstubin(VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_read_add),
.outervmstubin(VMS_L4D4PHI4X2n2_TE_L3D4PHI3X2_L4D4PHI4X2),
.number_in_innervmstubin(VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_number),
.read_add_innervmstubin(VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2_read_add),
.innervmstubin(VMS_L3D4PHI3X2n2_TE_L3D4PHI3X2_L4D4PHI4X2),
.stubpairout(TE_L3D4PHI3X2_L4D4PHI4X2_SP_L3D4PHI3X2_L4D4PHI4X2),
.valid_data(TE_L3D4PHI3X2_L4D4PHI4X2_SP_L3D4PHI3X2_L4D4PHI4X2_wr_en),
.start(VMS_L4D4PHI4X2n2_start),
.done(TE_L3D4PHI3X2_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI1X1_L6D3PHI1X1_phi.txt","TETable_TE_L5D3PHI1X1_L6D3PHI1X1_z.txt") TE_L5D3PHI1X1_L6D3PHI1X1(
.number_in_innervmstubin(VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_number),
.read_add_innervmstubin(VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_read_add),
.innervmstubin(VMS_L5D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1),
.number_in_outervmstubin(VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_number),
.read_add_outervmstubin(VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1_read_add),
.outervmstubin(VMS_L6D3PHI1X1n1_TE_L5D3PHI1X1_L6D3PHI1X1),
.stubpairout(TE_L5D3PHI1X1_L6D3PHI1X1_SP_L5D3PHI1X1_L6D3PHI1X1),
.valid_data(TE_L5D3PHI1X1_L6D3PHI1X1_SP_L5D3PHI1X1_L6D3PHI1X1_wr_en),
.start(VMS_L5D3PHI1X1n1_start),
.done(TE_L5D3PHI1X1_L6D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI1X1_L6D3PHI2X1_phi.txt","TETable_TE_L5D3PHI1X1_L6D3PHI2X1_z.txt") TE_L5D3PHI1X1_L6D3PHI2X1(
.number_in_innervmstubin(VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1_number),
.read_add_innervmstubin(VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1_read_add),
.innervmstubin(VMS_L5D3PHI1X1n2_TE_L5D3PHI1X1_L6D3PHI2X1),
.number_in_outervmstubin(VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1_number),
.read_add_outervmstubin(VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1_read_add),
.outervmstubin(VMS_L6D3PHI2X1n1_TE_L5D3PHI1X1_L6D3PHI2X1),
.stubpairout(TE_L5D3PHI1X1_L6D3PHI2X1_SP_L5D3PHI1X1_L6D3PHI2X1),
.valid_data(TE_L5D3PHI1X1_L6D3PHI2X1_SP_L5D3PHI1X1_L6D3PHI2X1_wr_en),
.start(VMS_L5D3PHI1X1n2_start),
.done(TE_L5D3PHI1X1_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI2X1_L6D3PHI2X1_phi.txt","TETable_TE_L5D3PHI2X1_L6D3PHI2X1_z.txt") TE_L5D3PHI2X1_L6D3PHI2X1(
.number_in_outervmstubin(VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1_number),
.read_add_outervmstubin(VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1_read_add),
.outervmstubin(VMS_L6D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI2X1),
.number_in_innervmstubin(VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1_number),
.read_add_innervmstubin(VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1_read_add),
.innervmstubin(VMS_L5D3PHI2X1n1_TE_L5D3PHI2X1_L6D3PHI2X1),
.stubpairout(TE_L5D3PHI2X1_L6D3PHI2X1_SP_L5D3PHI2X1_L6D3PHI2X1),
.valid_data(TE_L5D3PHI2X1_L6D3PHI2X1_SP_L5D3PHI2X1_L6D3PHI2X1_wr_en),
.start(VMS_L6D3PHI2X1n2_start),
.done(TE_L5D3PHI2X1_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI2X1_L6D3PHI3X1_phi.txt","TETable_TE_L5D3PHI2X1_L6D3PHI3X1_z.txt") TE_L5D3PHI2X1_L6D3PHI3X1(
.number_in_innervmstubin(VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1_number),
.read_add_innervmstubin(VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1_read_add),
.innervmstubin(VMS_L5D3PHI2X1n2_TE_L5D3PHI2X1_L6D3PHI3X1),
.number_in_outervmstubin(VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1_number),
.read_add_outervmstubin(VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1_read_add),
.outervmstubin(VMS_L6D3PHI3X1n1_TE_L5D3PHI2X1_L6D3PHI3X1),
.stubpairout(TE_L5D3PHI2X1_L6D3PHI3X1_SP_L5D3PHI2X1_L6D3PHI3X1),
.valid_data(TE_L5D3PHI2X1_L6D3PHI3X1_SP_L5D3PHI2X1_L6D3PHI3X1_wr_en),
.start(VMS_L5D3PHI2X1n2_start),
.done(TE_L5D3PHI2X1_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI3X1_L6D3PHI3X1_phi.txt","TETable_TE_L5D3PHI3X1_L6D3PHI3X1_z.txt") TE_L5D3PHI3X1_L6D3PHI3X1(
.number_in_outervmstubin(VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1_number),
.read_add_outervmstubin(VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1_read_add),
.outervmstubin(VMS_L6D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI3X1),
.number_in_innervmstubin(VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1_number),
.read_add_innervmstubin(VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1_read_add),
.innervmstubin(VMS_L5D3PHI3X1n1_TE_L5D3PHI3X1_L6D3PHI3X1),
.stubpairout(TE_L5D3PHI3X1_L6D3PHI3X1_SP_L5D3PHI3X1_L6D3PHI3X1),
.valid_data(TE_L5D3PHI3X1_L6D3PHI3X1_SP_L5D3PHI3X1_L6D3PHI3X1_wr_en),
.start(VMS_L6D3PHI3X1n2_start),
.done(TE_L5D3PHI3X1_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI3X1_L6D3PHI4X1_phi.txt","TETable_TE_L5D3PHI3X1_L6D3PHI4X1_z.txt") TE_L5D3PHI3X1_L6D3PHI4X1(
.number_in_innervmstubin(VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1_number),
.read_add_innervmstubin(VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1_read_add),
.innervmstubin(VMS_L5D3PHI3X1n2_TE_L5D3PHI3X1_L6D3PHI4X1),
.number_in_outervmstubin(VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1_number),
.read_add_outervmstubin(VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1_read_add),
.outervmstubin(VMS_L6D3PHI4X1n1_TE_L5D3PHI3X1_L6D3PHI4X1),
.stubpairout(TE_L5D3PHI3X1_L6D3PHI4X1_SP_L5D3PHI3X1_L6D3PHI4X1),
.valid_data(TE_L5D3PHI3X1_L6D3PHI4X1_SP_L5D3PHI3X1_L6D3PHI4X1_wr_en),
.start(VMS_L5D3PHI3X1n2_start),
.done(TE_L5D3PHI3X1_L6D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI1X1_L6D3PHI1X2_phi.txt","TETable_TE_L5D3PHI1X1_L6D3PHI1X2_z.txt") TE_L5D3PHI1X1_L6D3PHI1X2(
.number_in_innervmstubin(VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2_number),
.read_add_innervmstubin(VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2_read_add),
.innervmstubin(VMS_L5D3PHI1X1n3_TE_L5D3PHI1X1_L6D3PHI1X2),
.number_in_outervmstubin(VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2_number),
.read_add_outervmstubin(VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2_read_add),
.outervmstubin(VMS_L6D3PHI1X2n1_TE_L5D3PHI1X1_L6D3PHI1X2),
.stubpairout(TE_L5D3PHI1X1_L6D3PHI1X2_SP_L5D3PHI1X1_L6D3PHI1X2),
.valid_data(TE_L5D3PHI1X1_L6D3PHI1X2_SP_L5D3PHI1X1_L6D3PHI1X2_wr_en),
.start(VMS_L5D3PHI1X1n3_start),
.done(TE_L5D3PHI1X1_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI1X1_L6D3PHI2X2_phi.txt","TETable_TE_L5D3PHI1X1_L6D3PHI2X2_z.txt") TE_L5D3PHI1X1_L6D3PHI2X2(
.number_in_innervmstubin(VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2_number),
.read_add_innervmstubin(VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2_read_add),
.innervmstubin(VMS_L5D3PHI1X1n4_TE_L5D3PHI1X1_L6D3PHI2X2),
.number_in_outervmstubin(VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2_number),
.read_add_outervmstubin(VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2_read_add),
.outervmstubin(VMS_L6D3PHI2X2n1_TE_L5D3PHI1X1_L6D3PHI2X2),
.stubpairout(TE_L5D3PHI1X1_L6D3PHI2X2_SP_L5D3PHI1X1_L6D3PHI2X2),
.valid_data(TE_L5D3PHI1X1_L6D3PHI2X2_SP_L5D3PHI1X1_L6D3PHI2X2_wr_en),
.start(VMS_L5D3PHI1X1n4_start),
.done(TE_L5D3PHI1X1_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI2X1_L6D3PHI2X2_phi.txt","TETable_TE_L5D3PHI2X1_L6D3PHI2X2_z.txt") TE_L5D3PHI2X1_L6D3PHI2X2(
.number_in_innervmstubin(VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2_number),
.read_add_innervmstubin(VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2_read_add),
.innervmstubin(VMS_L5D3PHI2X1n3_TE_L5D3PHI2X1_L6D3PHI2X2),
.number_in_outervmstubin(VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2_number),
.read_add_outervmstubin(VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2_read_add),
.outervmstubin(VMS_L6D3PHI2X2n2_TE_L5D3PHI2X1_L6D3PHI2X2),
.stubpairout(TE_L5D3PHI2X1_L6D3PHI2X2_SP_L5D3PHI2X1_L6D3PHI2X2),
.valid_data(TE_L5D3PHI2X1_L6D3PHI2X2_SP_L5D3PHI2X1_L6D3PHI2X2_wr_en),
.start(VMS_L5D3PHI2X1n3_start),
.done(TE_L5D3PHI2X1_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI2X1_L6D3PHI3X2_phi.txt","TETable_TE_L5D3PHI2X1_L6D3PHI3X2_z.txt") TE_L5D3PHI2X1_L6D3PHI3X2(
.number_in_innervmstubin(VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2_number),
.read_add_innervmstubin(VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2_read_add),
.innervmstubin(VMS_L5D3PHI2X1n4_TE_L5D3PHI2X1_L6D3PHI3X2),
.number_in_outervmstubin(VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2_number),
.read_add_outervmstubin(VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2_read_add),
.outervmstubin(VMS_L6D3PHI3X2n1_TE_L5D3PHI2X1_L6D3PHI3X2),
.stubpairout(TE_L5D3PHI2X1_L6D3PHI3X2_SP_L5D3PHI2X1_L6D3PHI3X2),
.valid_data(TE_L5D3PHI2X1_L6D3PHI3X2_SP_L5D3PHI2X1_L6D3PHI3X2_wr_en),
.start(VMS_L5D3PHI2X1n4_start),
.done(TE_L5D3PHI2X1_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI3X1_L6D3PHI3X2_phi.txt","TETable_TE_L5D3PHI3X1_L6D3PHI3X2_z.txt") TE_L5D3PHI3X1_L6D3PHI3X2(
.number_in_innervmstubin(VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2_number),
.read_add_innervmstubin(VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2_read_add),
.innervmstubin(VMS_L5D3PHI3X1n3_TE_L5D3PHI3X1_L6D3PHI3X2),
.number_in_outervmstubin(VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2_number),
.read_add_outervmstubin(VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2_read_add),
.outervmstubin(VMS_L6D3PHI3X2n2_TE_L5D3PHI3X1_L6D3PHI3X2),
.stubpairout(TE_L5D3PHI3X1_L6D3PHI3X2_SP_L5D3PHI3X1_L6D3PHI3X2),
.valid_data(TE_L5D3PHI3X1_L6D3PHI3X2_SP_L5D3PHI3X1_L6D3PHI3X2_wr_en),
.start(VMS_L5D3PHI3X1n3_start),
.done(TE_L5D3PHI3X1_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI3X1_L6D3PHI4X2_phi.txt","TETable_TE_L5D3PHI3X1_L6D3PHI4X2_z.txt") TE_L5D3PHI3X1_L6D3PHI4X2(
.number_in_innervmstubin(VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2_number),
.read_add_innervmstubin(VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2_read_add),
.innervmstubin(VMS_L5D3PHI3X1n4_TE_L5D3PHI3X1_L6D3PHI4X2),
.number_in_outervmstubin(VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2_number),
.read_add_outervmstubin(VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2_read_add),
.outervmstubin(VMS_L6D3PHI4X2n1_TE_L5D3PHI3X1_L6D3PHI4X2),
.stubpairout(TE_L5D3PHI3X1_L6D3PHI4X2_SP_L5D3PHI3X1_L6D3PHI4X2),
.valid_data(TE_L5D3PHI3X1_L6D3PHI4X2_SP_L5D3PHI3X1_L6D3PHI4X2_wr_en),
.start(VMS_L5D3PHI3X1n4_start),
.done(TE_L5D3PHI3X1_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI1X2_L6D3PHI1X2_phi.txt","TETable_TE_L5D3PHI1X2_L6D3PHI1X2_z.txt") TE_L5D3PHI1X2_L6D3PHI1X2(
.number_in_outervmstubin(VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2_number),
.read_add_outervmstubin(VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2_read_add),
.outervmstubin(VMS_L6D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI1X2),
.number_in_innervmstubin(VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2_number),
.read_add_innervmstubin(VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2_read_add),
.innervmstubin(VMS_L5D3PHI1X2n1_TE_L5D3PHI1X2_L6D3PHI1X2),
.stubpairout(TE_L5D3PHI1X2_L6D3PHI1X2_SP_L5D3PHI1X2_L6D3PHI1X2),
.valid_data(TE_L5D3PHI1X2_L6D3PHI1X2_SP_L5D3PHI1X2_L6D3PHI1X2_wr_en),
.start(VMS_L6D3PHI1X2n2_start),
.done(TE_L5D3PHI1X2_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI1X2_L6D3PHI2X2_phi.txt","TETable_TE_L5D3PHI1X2_L6D3PHI2X2_z.txt") TE_L5D3PHI1X2_L6D3PHI2X2(
.number_in_outervmstubin(VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2_number),
.read_add_outervmstubin(VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2_read_add),
.outervmstubin(VMS_L6D3PHI2X2n3_TE_L5D3PHI1X2_L6D3PHI2X2),
.number_in_innervmstubin(VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2_number),
.read_add_innervmstubin(VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2_read_add),
.innervmstubin(VMS_L5D3PHI1X2n2_TE_L5D3PHI1X2_L6D3PHI2X2),
.stubpairout(TE_L5D3PHI1X2_L6D3PHI2X2_SP_L5D3PHI1X2_L6D3PHI2X2),
.valid_data(TE_L5D3PHI1X2_L6D3PHI2X2_SP_L5D3PHI1X2_L6D3PHI2X2_wr_en),
.start(VMS_L6D3PHI2X2n3_start),
.done(TE_L5D3PHI1X2_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI2X2_L6D3PHI2X2_phi.txt","TETable_TE_L5D3PHI2X2_L6D3PHI2X2_z.txt") TE_L5D3PHI2X2_L6D3PHI2X2(
.number_in_outervmstubin(VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2_number),
.read_add_outervmstubin(VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2_read_add),
.outervmstubin(VMS_L6D3PHI2X2n4_TE_L5D3PHI2X2_L6D3PHI2X2),
.number_in_innervmstubin(VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2_number),
.read_add_innervmstubin(VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2_read_add),
.innervmstubin(VMS_L5D3PHI2X2n1_TE_L5D3PHI2X2_L6D3PHI2X2),
.stubpairout(TE_L5D3PHI2X2_L6D3PHI2X2_SP_L5D3PHI2X2_L6D3PHI2X2),
.valid_data(TE_L5D3PHI2X2_L6D3PHI2X2_SP_L5D3PHI2X2_L6D3PHI2X2_wr_en),
.start(VMS_L6D3PHI2X2n4_start),
.done(TE_L5D3PHI2X2_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI2X2_L6D3PHI3X2_phi.txt","TETable_TE_L5D3PHI2X2_L6D3PHI3X2_z.txt") TE_L5D3PHI2X2_L6D3PHI3X2(
.number_in_outervmstubin(VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2_number),
.read_add_outervmstubin(VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2_read_add),
.outervmstubin(VMS_L6D3PHI3X2n3_TE_L5D3PHI2X2_L6D3PHI3X2),
.number_in_innervmstubin(VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2_number),
.read_add_innervmstubin(VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2_read_add),
.innervmstubin(VMS_L5D3PHI2X2n2_TE_L5D3PHI2X2_L6D3PHI3X2),
.stubpairout(TE_L5D3PHI2X2_L6D3PHI3X2_SP_L5D3PHI2X2_L6D3PHI3X2),
.valid_data(TE_L5D3PHI2X2_L6D3PHI3X2_SP_L5D3PHI2X2_L6D3PHI3X2_wr_en),
.start(VMS_L6D3PHI3X2n3_start),
.done(TE_L5D3PHI2X2_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI3X2_L6D3PHI3X2_phi.txt","TETable_TE_L5D3PHI3X2_L6D3PHI3X2_z.txt") TE_L5D3PHI3X2_L6D3PHI3X2(
.number_in_outervmstubin(VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2_number),
.read_add_outervmstubin(VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2_read_add),
.outervmstubin(VMS_L6D3PHI3X2n4_TE_L5D3PHI3X2_L6D3PHI3X2),
.number_in_innervmstubin(VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2_number),
.read_add_innervmstubin(VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2_read_add),
.innervmstubin(VMS_L5D3PHI3X2n1_TE_L5D3PHI3X2_L6D3PHI3X2),
.stubpairout(TE_L5D3PHI3X2_L6D3PHI3X2_SP_L5D3PHI3X2_L6D3PHI3X2),
.valid_data(TE_L5D3PHI3X2_L6D3PHI3X2_SP_L5D3PHI3X2_L6D3PHI3X2_wr_en),
.start(VMS_L6D3PHI3X2n4_start),
.done(TE_L5D3PHI3X2_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI3X2_L6D3PHI4X2_phi.txt","TETable_TE_L5D3PHI3X2_L6D3PHI4X2_z.txt") TE_L5D3PHI3X2_L6D3PHI4X2(
.number_in_outervmstubin(VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_number),
.read_add_outervmstubin(VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_read_add),
.outervmstubin(VMS_L6D3PHI4X2n2_TE_L5D3PHI3X2_L6D3PHI4X2),
.number_in_innervmstubin(VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_number),
.read_add_innervmstubin(VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2_read_add),
.innervmstubin(VMS_L5D3PHI3X2n2_TE_L5D3PHI3X2_L6D3PHI4X2),
.stubpairout(TE_L5D3PHI3X2_L6D3PHI4X2_SP_L5D3PHI3X2_L6D3PHI4X2),
.valid_data(TE_L5D3PHI3X2_L6D3PHI4X2_SP_L5D3PHI3X2_L6D3PHI4X2_wr_en),
.start(VMS_L6D3PHI4X2n2_start),
.done(TE_L5D3PHI3X2_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI1X2_L6D4PHI1X1_phi.txt","TETable_TE_L5D3PHI1X2_L6D4PHI1X1_z.txt") TE_L5D3PHI1X2_L6D4PHI1X1(
.number_in_innervmstubin(VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1_number),
.read_add_innervmstubin(VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1_read_add),
.innervmstubin(VMS_L5D3PHI1X2n3_TE_L5D3PHI1X2_L6D4PHI1X1),
.number_in_outervmstubin(VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1_number),
.read_add_outervmstubin(VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1_read_add),
.outervmstubin(VMS_L6D4PHI1X1n1_TE_L5D3PHI1X2_L6D4PHI1X1),
.stubpairout(TE_L5D3PHI1X2_L6D4PHI1X1_SP_L5D3PHI1X2_L6D4PHI1X1),
.valid_data(TE_L5D3PHI1X2_L6D4PHI1X1_SP_L5D3PHI1X2_L6D4PHI1X1_wr_en),
.start(VMS_L5D3PHI1X2n3_start),
.done(TE_L5D3PHI1X2_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI1X2_L6D4PHI2X1_phi.txt","TETable_TE_L5D3PHI1X2_L6D4PHI2X1_z.txt") TE_L5D3PHI1X2_L6D4PHI2X1(
.number_in_innervmstubin(VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1_number),
.read_add_innervmstubin(VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1_read_add),
.innervmstubin(VMS_L5D3PHI1X2n4_TE_L5D3PHI1X2_L6D4PHI2X1),
.number_in_outervmstubin(VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1_number),
.read_add_outervmstubin(VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1_read_add),
.outervmstubin(VMS_L6D4PHI2X1n1_TE_L5D3PHI1X2_L6D4PHI2X1),
.stubpairout(TE_L5D3PHI1X2_L6D4PHI2X1_SP_L5D3PHI1X2_L6D4PHI2X1),
.valid_data(TE_L5D3PHI1X2_L6D4PHI2X1_SP_L5D3PHI1X2_L6D4PHI2X1_wr_en),
.start(VMS_L5D3PHI1X2n4_start),
.done(TE_L5D3PHI1X2_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI2X2_L6D4PHI2X1_phi.txt","TETable_TE_L5D3PHI2X2_L6D4PHI2X1_z.txt") TE_L5D3PHI2X2_L6D4PHI2X1(
.number_in_innervmstubin(VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1_number),
.read_add_innervmstubin(VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1_read_add),
.innervmstubin(VMS_L5D3PHI2X2n3_TE_L5D3PHI2X2_L6D4PHI2X1),
.number_in_outervmstubin(VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1_number),
.read_add_outervmstubin(VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1_read_add),
.outervmstubin(VMS_L6D4PHI2X1n2_TE_L5D3PHI2X2_L6D4PHI2X1),
.stubpairout(TE_L5D3PHI2X2_L6D4PHI2X1_SP_L5D3PHI2X2_L6D4PHI2X1),
.valid_data(TE_L5D3PHI2X2_L6D4PHI2X1_SP_L5D3PHI2X2_L6D4PHI2X1_wr_en),
.start(VMS_L5D3PHI2X2n3_start),
.done(TE_L5D3PHI2X2_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI2X2_L6D4PHI3X1_phi.txt","TETable_TE_L5D3PHI2X2_L6D4PHI3X1_z.txt") TE_L5D3PHI2X2_L6D4PHI3X1(
.number_in_innervmstubin(VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1_number),
.read_add_innervmstubin(VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1_read_add),
.innervmstubin(VMS_L5D3PHI2X2n4_TE_L5D3PHI2X2_L6D4PHI3X1),
.number_in_outervmstubin(VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1_number),
.read_add_outervmstubin(VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1_read_add),
.outervmstubin(VMS_L6D4PHI3X1n1_TE_L5D3PHI2X2_L6D4PHI3X1),
.stubpairout(TE_L5D3PHI2X2_L6D4PHI3X1_SP_L5D3PHI2X2_L6D4PHI3X1),
.valid_data(TE_L5D3PHI2X2_L6D4PHI3X1_SP_L5D3PHI2X2_L6D4PHI3X1_wr_en),
.start(VMS_L5D3PHI2X2n4_start),
.done(TE_L5D3PHI2X2_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI3X2_L6D4PHI3X1_phi.txt","TETable_TE_L5D3PHI3X2_L6D4PHI3X1_z.txt") TE_L5D3PHI3X2_L6D4PHI3X1(
.number_in_innervmstubin(VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1_number),
.read_add_innervmstubin(VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1_read_add),
.innervmstubin(VMS_L5D3PHI3X2n3_TE_L5D3PHI3X2_L6D4PHI3X1),
.number_in_outervmstubin(VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1_number),
.read_add_outervmstubin(VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1_read_add),
.outervmstubin(VMS_L6D4PHI3X1n2_TE_L5D3PHI3X2_L6D4PHI3X1),
.stubpairout(TE_L5D3PHI3X2_L6D4PHI3X1_SP_L5D3PHI3X2_L6D4PHI3X1),
.valid_data(TE_L5D3PHI3X2_L6D4PHI3X1_SP_L5D3PHI3X2_L6D4PHI3X1_wr_en),
.start(VMS_L5D3PHI3X2n3_start),
.done(TE_L5D3PHI3X2_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D3PHI3X2_L6D4PHI4X1_phi.txt","TETable_TE_L5D3PHI3X2_L6D4PHI4X1_z.txt") TE_L5D3PHI3X2_L6D4PHI4X1(
.number_in_innervmstubin(VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1_number),
.read_add_innervmstubin(VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1_read_add),
.innervmstubin(VMS_L5D3PHI3X2n4_TE_L5D3PHI3X2_L6D4PHI4X1),
.number_in_outervmstubin(VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1_number),
.read_add_outervmstubin(VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1_read_add),
.outervmstubin(VMS_L6D4PHI4X1n1_TE_L5D3PHI3X2_L6D4PHI4X1),
.stubpairout(TE_L5D3PHI3X2_L6D4PHI4X1_SP_L5D3PHI3X2_L6D4PHI4X1),
.valid_data(TE_L5D3PHI3X2_L6D4PHI4X1_SP_L5D3PHI3X2_L6D4PHI4X1_wr_en),
.start(VMS_L5D3PHI3X2n4_start),
.done(TE_L5D3PHI3X2_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI1X1_L6D4PHI1X1_phi.txt","TETable_TE_L5D4PHI1X1_L6D4PHI1X1_z.txt") TE_L5D4PHI1X1_L6D4PHI1X1(
.number_in_outervmstubin(VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1_number),
.read_add_outervmstubin(VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1_read_add),
.outervmstubin(VMS_L6D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI1X1),
.number_in_innervmstubin(VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1_number),
.read_add_innervmstubin(VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1_read_add),
.innervmstubin(VMS_L5D4PHI1X1n1_TE_L5D4PHI1X1_L6D4PHI1X1),
.stubpairout(TE_L5D4PHI1X1_L6D4PHI1X1_SP_L5D4PHI1X1_L6D4PHI1X1),
.valid_data(TE_L5D4PHI1X1_L6D4PHI1X1_SP_L5D4PHI1X1_L6D4PHI1X1_wr_en),
.start(VMS_L6D4PHI1X1n2_start),
.done(TE_L5D4PHI1X1_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI1X1_L6D4PHI2X1_phi.txt","TETable_TE_L5D4PHI1X1_L6D4PHI2X1_z.txt") TE_L5D4PHI1X1_L6D4PHI2X1(
.number_in_outervmstubin(VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1_number),
.read_add_outervmstubin(VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1_read_add),
.outervmstubin(VMS_L6D4PHI2X1n3_TE_L5D4PHI1X1_L6D4PHI2X1),
.number_in_innervmstubin(VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1_number),
.read_add_innervmstubin(VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1_read_add),
.innervmstubin(VMS_L5D4PHI1X1n2_TE_L5D4PHI1X1_L6D4PHI2X1),
.stubpairout(TE_L5D4PHI1X1_L6D4PHI2X1_SP_L5D4PHI1X1_L6D4PHI2X1),
.valid_data(TE_L5D4PHI1X1_L6D4PHI2X1_SP_L5D4PHI1X1_L6D4PHI2X1_wr_en),
.start(VMS_L6D4PHI2X1n3_start),
.done(TE_L5D4PHI1X1_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI2X1_L6D4PHI2X1_phi.txt","TETable_TE_L5D4PHI2X1_L6D4PHI2X1_z.txt") TE_L5D4PHI2X1_L6D4PHI2X1(
.number_in_outervmstubin(VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1_number),
.read_add_outervmstubin(VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1_read_add),
.outervmstubin(VMS_L6D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI2X1),
.number_in_innervmstubin(VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1_number),
.read_add_innervmstubin(VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1_read_add),
.innervmstubin(VMS_L5D4PHI2X1n1_TE_L5D4PHI2X1_L6D4PHI2X1),
.stubpairout(TE_L5D4PHI2X1_L6D4PHI2X1_SP_L5D4PHI2X1_L6D4PHI2X1),
.valid_data(TE_L5D4PHI2X1_L6D4PHI2X1_SP_L5D4PHI2X1_L6D4PHI2X1_wr_en),
.start(VMS_L6D4PHI2X1n4_start),
.done(TE_L5D4PHI2X1_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI2X1_L6D4PHI3X1_phi.txt","TETable_TE_L5D4PHI2X1_L6D4PHI3X1_z.txt") TE_L5D4PHI2X1_L6D4PHI3X1(
.number_in_outervmstubin(VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1_number),
.read_add_outervmstubin(VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1_read_add),
.outervmstubin(VMS_L6D4PHI3X1n3_TE_L5D4PHI2X1_L6D4PHI3X1),
.number_in_innervmstubin(VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1_number),
.read_add_innervmstubin(VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1_read_add),
.innervmstubin(VMS_L5D4PHI2X1n2_TE_L5D4PHI2X1_L6D4PHI3X1),
.stubpairout(TE_L5D4PHI2X1_L6D4PHI3X1_SP_L5D4PHI2X1_L6D4PHI3X1),
.valid_data(TE_L5D4PHI2X1_L6D4PHI3X1_SP_L5D4PHI2X1_L6D4PHI3X1_wr_en),
.start(VMS_L6D4PHI3X1n3_start),
.done(TE_L5D4PHI2X1_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI3X1_L6D4PHI3X1_phi.txt","TETable_TE_L5D4PHI3X1_L6D4PHI3X1_z.txt") TE_L5D4PHI3X1_L6D4PHI3X1(
.number_in_outervmstubin(VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1_number),
.read_add_outervmstubin(VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1_read_add),
.outervmstubin(VMS_L6D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI3X1),
.number_in_innervmstubin(VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1_number),
.read_add_innervmstubin(VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1_read_add),
.innervmstubin(VMS_L5D4PHI3X1n1_TE_L5D4PHI3X1_L6D4PHI3X1),
.stubpairout(TE_L5D4PHI3X1_L6D4PHI3X1_SP_L5D4PHI3X1_L6D4PHI3X1),
.valid_data(TE_L5D4PHI3X1_L6D4PHI3X1_SP_L5D4PHI3X1_L6D4PHI3X1_wr_en),
.start(VMS_L6D4PHI3X1n4_start),
.done(TE_L5D4PHI3X1_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI3X1_L6D4PHI4X1_phi.txt","TETable_TE_L5D4PHI3X1_L6D4PHI4X1_z.txt") TE_L5D4PHI3X1_L6D4PHI4X1(
.number_in_outervmstubin(VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_number),
.read_add_outervmstubin(VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_read_add),
.outervmstubin(VMS_L6D4PHI4X1n2_TE_L5D4PHI3X1_L6D4PHI4X1),
.number_in_innervmstubin(VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_number),
.read_add_innervmstubin(VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1_read_add),
.innervmstubin(VMS_L5D4PHI3X1n2_TE_L5D4PHI3X1_L6D4PHI4X1),
.stubpairout(TE_L5D4PHI3X1_L6D4PHI4X1_SP_L5D4PHI3X1_L6D4PHI4X1),
.valid_data(TE_L5D4PHI3X1_L6D4PHI4X1_SP_L5D4PHI3X1_L6D4PHI4X1_wr_en),
.start(VMS_L6D4PHI4X1n2_start),
.done(TE_L5D4PHI3X1_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI1X1_L6D4PHI1X2_phi.txt","TETable_TE_L5D4PHI1X1_L6D4PHI1X2_z.txt") TE_L5D4PHI1X1_L6D4PHI1X2(
.number_in_innervmstubin(VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2_number),
.read_add_innervmstubin(VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2_read_add),
.innervmstubin(VMS_L5D4PHI1X1n3_TE_L5D4PHI1X1_L6D4PHI1X2),
.number_in_outervmstubin(VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2_number),
.read_add_outervmstubin(VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2_read_add),
.outervmstubin(VMS_L6D4PHI1X2n1_TE_L5D4PHI1X1_L6D4PHI1X2),
.stubpairout(TE_L5D4PHI1X1_L6D4PHI1X2_SP_L5D4PHI1X1_L6D4PHI1X2),
.valid_data(TE_L5D4PHI1X1_L6D4PHI1X2_SP_L5D4PHI1X1_L6D4PHI1X2_wr_en),
.start(VMS_L5D4PHI1X1n3_start),
.done(TE_L5D4PHI1X1_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI1X1_L6D4PHI2X2_phi.txt","TETable_TE_L5D4PHI1X1_L6D4PHI2X2_z.txt") TE_L5D4PHI1X1_L6D4PHI2X2(
.number_in_innervmstubin(VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2_number),
.read_add_innervmstubin(VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2_read_add),
.innervmstubin(VMS_L5D4PHI1X1n4_TE_L5D4PHI1X1_L6D4PHI2X2),
.number_in_outervmstubin(VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2_number),
.read_add_outervmstubin(VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2_read_add),
.outervmstubin(VMS_L6D4PHI2X2n1_TE_L5D4PHI1X1_L6D4PHI2X2),
.stubpairout(TE_L5D4PHI1X1_L6D4PHI2X2_SP_L5D4PHI1X1_L6D4PHI2X2),
.valid_data(TE_L5D4PHI1X1_L6D4PHI2X2_SP_L5D4PHI1X1_L6D4PHI2X2_wr_en),
.start(VMS_L5D4PHI1X1n4_start),
.done(TE_L5D4PHI1X1_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI2X1_L6D4PHI2X2_phi.txt","TETable_TE_L5D4PHI2X1_L6D4PHI2X2_z.txt") TE_L5D4PHI2X1_L6D4PHI2X2(
.number_in_innervmstubin(VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2_number),
.read_add_innervmstubin(VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2_read_add),
.innervmstubin(VMS_L5D4PHI2X1n3_TE_L5D4PHI2X1_L6D4PHI2X2),
.number_in_outervmstubin(VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2_number),
.read_add_outervmstubin(VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2_read_add),
.outervmstubin(VMS_L6D4PHI2X2n2_TE_L5D4PHI2X1_L6D4PHI2X2),
.stubpairout(TE_L5D4PHI2X1_L6D4PHI2X2_SP_L5D4PHI2X1_L6D4PHI2X2),
.valid_data(TE_L5D4PHI2X1_L6D4PHI2X2_SP_L5D4PHI2X1_L6D4PHI2X2_wr_en),
.start(VMS_L5D4PHI2X1n3_start),
.done(TE_L5D4PHI2X1_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI2X1_L6D4PHI3X2_phi.txt","TETable_TE_L5D4PHI2X1_L6D4PHI3X2_z.txt") TE_L5D4PHI2X1_L6D4PHI3X2(
.number_in_innervmstubin(VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2_number),
.read_add_innervmstubin(VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2_read_add),
.innervmstubin(VMS_L5D4PHI2X1n4_TE_L5D4PHI2X1_L6D4PHI3X2),
.number_in_outervmstubin(VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2_number),
.read_add_outervmstubin(VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2_read_add),
.outervmstubin(VMS_L6D4PHI3X2n1_TE_L5D4PHI2X1_L6D4PHI3X2),
.stubpairout(TE_L5D4PHI2X1_L6D4PHI3X2_SP_L5D4PHI2X1_L6D4PHI3X2),
.valid_data(TE_L5D4PHI2X1_L6D4PHI3X2_SP_L5D4PHI2X1_L6D4PHI3X2_wr_en),
.start(VMS_L5D4PHI2X1n4_start),
.done(TE_L5D4PHI2X1_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI3X1_L6D4PHI3X2_phi.txt","TETable_TE_L5D4PHI3X1_L6D4PHI3X2_z.txt") TE_L5D4PHI3X1_L6D4PHI3X2(
.number_in_innervmstubin(VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2_number),
.read_add_innervmstubin(VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2_read_add),
.innervmstubin(VMS_L5D4PHI3X1n3_TE_L5D4PHI3X1_L6D4PHI3X2),
.number_in_outervmstubin(VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2_number),
.read_add_outervmstubin(VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2_read_add),
.outervmstubin(VMS_L6D4PHI3X2n2_TE_L5D4PHI3X1_L6D4PHI3X2),
.stubpairout(TE_L5D4PHI3X1_L6D4PHI3X2_SP_L5D4PHI3X1_L6D4PHI3X2),
.valid_data(TE_L5D4PHI3X1_L6D4PHI3X2_SP_L5D4PHI3X1_L6D4PHI3X2_wr_en),
.start(VMS_L5D4PHI3X1n3_start),
.done(TE_L5D4PHI3X1_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI3X1_L6D4PHI4X2_phi.txt","TETable_TE_L5D4PHI3X1_L6D4PHI4X2_z.txt") TE_L5D4PHI3X1_L6D4PHI4X2(
.number_in_innervmstubin(VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2_number),
.read_add_innervmstubin(VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2_read_add),
.innervmstubin(VMS_L5D4PHI3X1n4_TE_L5D4PHI3X1_L6D4PHI4X2),
.number_in_outervmstubin(VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2_number),
.read_add_outervmstubin(VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2_read_add),
.outervmstubin(VMS_L6D4PHI4X2n1_TE_L5D4PHI3X1_L6D4PHI4X2),
.stubpairout(TE_L5D4PHI3X1_L6D4PHI4X2_SP_L5D4PHI3X1_L6D4PHI4X2),
.valid_data(TE_L5D4PHI3X1_L6D4PHI4X2_SP_L5D4PHI3X1_L6D4PHI4X2_wr_en),
.start(VMS_L5D4PHI3X1n4_start),
.done(TE_L5D4PHI3X1_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI1X2_L6D4PHI1X2_phi.txt","TETable_TE_L5D4PHI1X2_L6D4PHI1X2_z.txt") TE_L5D4PHI1X2_L6D4PHI1X2(
.number_in_outervmstubin(VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2_number),
.read_add_outervmstubin(VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2_read_add),
.outervmstubin(VMS_L6D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI1X2),
.number_in_innervmstubin(VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2_number),
.read_add_innervmstubin(VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2_read_add),
.innervmstubin(VMS_L5D4PHI1X2n1_TE_L5D4PHI1X2_L6D4PHI1X2),
.stubpairout(TE_L5D4PHI1X2_L6D4PHI1X2_SP_L5D4PHI1X2_L6D4PHI1X2),
.valid_data(TE_L5D4PHI1X2_L6D4PHI1X2_SP_L5D4PHI1X2_L6D4PHI1X2_wr_en),
.start(VMS_L6D4PHI1X2n2_start),
.done(TE_L5D4PHI1X2_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI1X2_L6D4PHI2X2_phi.txt","TETable_TE_L5D4PHI1X2_L6D4PHI2X2_z.txt") TE_L5D4PHI1X2_L6D4PHI2X2(
.number_in_outervmstubin(VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2_number),
.read_add_outervmstubin(VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2_read_add),
.outervmstubin(VMS_L6D4PHI2X2n3_TE_L5D4PHI1X2_L6D4PHI2X2),
.number_in_innervmstubin(VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2_number),
.read_add_innervmstubin(VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2_read_add),
.innervmstubin(VMS_L5D4PHI1X2n2_TE_L5D4PHI1X2_L6D4PHI2X2),
.stubpairout(TE_L5D4PHI1X2_L6D4PHI2X2_SP_L5D4PHI1X2_L6D4PHI2X2),
.valid_data(TE_L5D4PHI1X2_L6D4PHI2X2_SP_L5D4PHI1X2_L6D4PHI2X2_wr_en),
.start(VMS_L6D4PHI2X2n3_start),
.done(TE_L5D4PHI1X2_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI2X2_L6D4PHI2X2_phi.txt","TETable_TE_L5D4PHI2X2_L6D4PHI2X2_z.txt") TE_L5D4PHI2X2_L6D4PHI2X2(
.number_in_outervmstubin(VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2_number),
.read_add_outervmstubin(VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2_read_add),
.outervmstubin(VMS_L6D4PHI2X2n4_TE_L5D4PHI2X2_L6D4PHI2X2),
.number_in_innervmstubin(VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2_number),
.read_add_innervmstubin(VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2_read_add),
.innervmstubin(VMS_L5D4PHI2X2n1_TE_L5D4PHI2X2_L6D4PHI2X2),
.stubpairout(TE_L5D4PHI2X2_L6D4PHI2X2_SP_L5D4PHI2X2_L6D4PHI2X2),
.valid_data(TE_L5D4PHI2X2_L6D4PHI2X2_SP_L5D4PHI2X2_L6D4PHI2X2_wr_en),
.start(VMS_L6D4PHI2X2n4_start),
.done(TE_L5D4PHI2X2_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI2X2_L6D4PHI3X2_phi.txt","TETable_TE_L5D4PHI2X2_L6D4PHI3X2_z.txt") TE_L5D4PHI2X2_L6D4PHI3X2(
.number_in_outervmstubin(VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2_number),
.read_add_outervmstubin(VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2_read_add),
.outervmstubin(VMS_L6D4PHI3X2n3_TE_L5D4PHI2X2_L6D4PHI3X2),
.number_in_innervmstubin(VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2_number),
.read_add_innervmstubin(VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2_read_add),
.innervmstubin(VMS_L5D4PHI2X2n2_TE_L5D4PHI2X2_L6D4PHI3X2),
.stubpairout(TE_L5D4PHI2X2_L6D4PHI3X2_SP_L5D4PHI2X2_L6D4PHI3X2),
.valid_data(TE_L5D4PHI2X2_L6D4PHI3X2_SP_L5D4PHI2X2_L6D4PHI3X2_wr_en),
.start(VMS_L6D4PHI3X2n3_start),
.done(TE_L5D4PHI2X2_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI3X2_L6D4PHI3X2_phi.txt","TETable_TE_L5D4PHI3X2_L6D4PHI3X2_z.txt") TE_L5D4PHI3X2_L6D4PHI3X2(
.number_in_outervmstubin(VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2_number),
.read_add_outervmstubin(VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2_read_add),
.outervmstubin(VMS_L6D4PHI3X2n4_TE_L5D4PHI3X2_L6D4PHI3X2),
.number_in_innervmstubin(VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2_number),
.read_add_innervmstubin(VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2_read_add),
.innervmstubin(VMS_L5D4PHI3X2n1_TE_L5D4PHI3X2_L6D4PHI3X2),
.stubpairout(TE_L5D4PHI3X2_L6D4PHI3X2_SP_L5D4PHI3X2_L6D4PHI3X2),
.valid_data(TE_L5D4PHI3X2_L6D4PHI3X2_SP_L5D4PHI3X2_L6D4PHI3X2_wr_en),
.start(VMS_L6D4PHI3X2n4_start),
.done(TE_L5D4PHI3X2_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletEngine #("TETable_TE_L5D4PHI3X2_L6D4PHI4X2_phi.txt","TETable_TE_L5D4PHI3X2_L6D4PHI4X2_z.txt") TE_L5D4PHI3X2_L6D4PHI4X2(
.number_in_outervmstubin(VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_number),
.read_add_outervmstubin(VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_read_add),
.outervmstubin(VMS_L6D4PHI4X2n2_TE_L5D4PHI3X2_L6D4PHI4X2),
.number_in_innervmstubin(VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_number),
.read_add_innervmstubin(VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2_read_add),
.innervmstubin(VMS_L5D4PHI3X2n2_TE_L5D4PHI3X2_L6D4PHI4X2),
.stubpairout(TE_L5D4PHI3X2_L6D4PHI4X2_SP_L5D4PHI3X2_L6D4PHI4X2),
.valid_data(TE_L5D4PHI3X2_L6D4PHI4X2_SP_L5D4PHI3X2_L6D4PHI4X2_wr_en),
.start(VMS_L6D4PHI4X2n2_start),
.done(TE_L5D4PHI3X2_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L1D3L2D3.dat"),.R1MEAN(`TC_L1L2_krA),.R2MEAN(`TC_L1L2_krB),.TC_index(4'b0000),.IsInner1(1'b1),.IsInner2(1'b1)) TC_L1D3L2D3(
.number_in_stubpair1in(SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3_number),
.read_add_stubpair1in(SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3_read_add),
.stubpair1in(SP_L1D3PHI1X1_L2D3PHI1X1_TC_L1D3L2D3),
.number_in_stubpair2in(SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3_number),
.read_add_stubpair2in(SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3_read_add),
.stubpair2in(SP_L1D3PHI1X1_L2D3PHI2X1_TC_L1D3L2D3),
.number_in_stubpair3in(SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3_number),
.read_add_stubpair3in(SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3_read_add),
.stubpair3in(SP_L1D3PHI2X1_L2D3PHI2X1_TC_L1D3L2D3),
.number_in_stubpair4in(SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3_number),
.read_add_stubpair4in(SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3_read_add),
.stubpair4in(SP_L1D3PHI2X1_L2D3PHI3X1_TC_L1D3L2D3),
.number_in_stubpair5in(SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3_number),
.read_add_stubpair5in(SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3_read_add),
.stubpair5in(SP_L1D3PHI3X1_L2D3PHI3X1_TC_L1D3L2D3),
.number_in_stubpair6in(SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3_number),
.read_add_stubpair6in(SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3_read_add),
.stubpair6in(SP_L1D3PHI3X1_L2D3PHI4X1_TC_L1D3L2D3),
.number_in_stubpair7in(SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3_number),
.read_add_stubpair7in(SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3_read_add),
.stubpair7in(SP_L1D3PHI1X1_L2D3PHI1X2_TC_L1D3L2D3),
.number_in_stubpair8in(SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3_number),
.read_add_stubpair8in(SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3_read_add),
.stubpair8in(SP_L1D3PHI1X1_L2D3PHI2X2_TC_L1D3L2D3),
.number_in_stubpair9in(SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3_number),
.read_add_stubpair9in(SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3_read_add),
.stubpair9in(SP_L1D3PHI2X1_L2D3PHI2X2_TC_L1D3L2D3),
.number_in_stubpair10in(SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3_number),
.read_add_stubpair10in(SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3_read_add),
.stubpair10in(SP_L1D3PHI2X1_L2D3PHI3X2_TC_L1D3L2D3),
.number_in_stubpair11in(SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3_number),
.read_add_stubpair11in(SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3_read_add),
.stubpair11in(SP_L1D3PHI3X1_L2D3PHI3X2_TC_L1D3L2D3),
.number_in_stubpair12in(SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3_number),
.read_add_stubpair12in(SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3_read_add),
.stubpair12in(SP_L1D3PHI3X1_L2D3PHI4X2_TC_L1D3L2D3),
.number_in_stubpair13in(SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3_number),
.read_add_stubpair13in(SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3_read_add),
.stubpair13in(SP_L1D3PHI1X2_L2D3PHI1X2_TC_L1D3L2D3),
.number_in_stubpair14in(SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3_number),
.read_add_stubpair14in(SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3_read_add),
.stubpair14in(SP_L1D3PHI1X2_L2D3PHI2X2_TC_L1D3L2D3),
.number_in_stubpair15in(SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3_number),
.read_add_stubpair15in(SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3_read_add),
.stubpair15in(SP_L1D3PHI2X2_L2D3PHI2X2_TC_L1D3L2D3),
.number_in_stubpair16in(SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3_number),
.read_add_stubpair16in(SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3_read_add),
.stubpair16in(SP_L1D3PHI2X2_L2D3PHI3X2_TC_L1D3L2D3),
.number_in_stubpair17in(SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3_number),
.read_add_stubpair17in(SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3_read_add),
.stubpair17in(SP_L1D3PHI3X2_L2D3PHI3X2_TC_L1D3L2D3),
.number_in_stubpair18in(SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3_number),
.read_add_stubpair18in(SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3_read_add),
.stubpair18in(SP_L1D3PHI3X2_L2D3PHI4X2_TC_L1D3L2D3),
.read_add_outerallstubin(AS_L2D3n1_TC_L1D3L2D3_read_add),
.outerallstubin(AS_L2D3n1_TC_L1D3L2D3),
.read_add_innerallstubin(AS_L1D3n1_TC_L1D3L2D3_read_add),
.innerallstubin(AS_L1D3n1_TC_L1D3L2D3),
.projoutToPlus_L3(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3),
.projoutToPlus_L4(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4),
.projoutToPlus_L5(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5),
.projoutToPlus_L6(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6),
.projoutToMinus_L3(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3),
.projoutToMinus_L4(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4),
.projoutToMinus_L5(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5),
.projoutToMinus_L6(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6),
.projout_L3D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3),
.projout_L4D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3),
.projout_L5D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3),
.projout_L6D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3),
.projout_L3D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4),
.projout_L4D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4),
.projout_L5D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4),
.projout_L6D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4),
.trackpar(TC_L1D3L2D3_TPAR_L1D3L2D3),
.valid_projoutToPlus_L3(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L3_wr_en),
.valid_projoutToPlus_L4(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L4_wr_en),
.valid_projoutToPlus_L5(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L5_wr_en),
.valid_projoutToPlus_L6(TC_L1D3L2D3_TPROJ_ToPlus_L1D3L2D3_L6_wr_en),
.valid_projoutToMinus_L3(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L3_wr_en),
.valid_projoutToMinus_L4(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L4_wr_en),
.valid_projoutToMinus_L5(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L5_wr_en),
.valid_projoutToMinus_L6(TC_L1D3L2D3_TPROJ_ToMinus_L1D3L2D3_L6_wr_en),
.valid_projout_L3D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D3_wr_en),
.valid_projout_L4D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D3_wr_en),
.valid_projout_L5D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D3_wr_en),
.valid_projout_L6D3(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D3_wr_en),
.valid_projout_L3D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L3D4_wr_en),
.valid_projout_L4D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L4D4_wr_en),
.valid_projout_L5D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L5D4_wr_en),
.valid_projout_L6D4(TC_L1D3L2D3_TPROJ_L1D3L2D3_L6D4_wr_en),
.valid_trackpar(TC_L1D3L2D3_TPAR_L1D3L2D3_wr_en),
.done_proj(TC_L1D3L2D3_proj_start),
.start(SP_L1D3PHI1X1_L2D3PHI1X1_start),
.done(TC_L1D3L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L1D3L2D3.dat"),.R1MEAN(`TC_L1L2_krA),.R2MEAN(`TC_L1L2_krB),.TC_index(4'b0001),.IsInner1(1'b1),.IsInner2(1'b1)) TC_L1D3L2D4(
.number_in_stubpair1in(SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4_number),
.read_add_stubpair1in(SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4_read_add),
.stubpair1in(SP_L1D3PHI1X1_L2D4PHI1X1_TC_L1D3L2D4),
.number_in_stubpair2in(SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4_number),
.read_add_stubpair2in(SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4_read_add),
.stubpair2in(SP_L1D3PHI1X1_L2D4PHI2X1_TC_L1D3L2D4),
.number_in_stubpair3in(SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4_number),
.read_add_stubpair3in(SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4_read_add),
.stubpair3in(SP_L1D3PHI2X1_L2D4PHI2X1_TC_L1D3L2D4),
.number_in_stubpair4in(SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4_number),
.read_add_stubpair4in(SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4_read_add),
.stubpair4in(SP_L1D3PHI2X1_L2D4PHI3X1_TC_L1D3L2D4),
.number_in_stubpair5in(SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4_number),
.read_add_stubpair5in(SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4_read_add),
.stubpair5in(SP_L1D3PHI3X1_L2D4PHI3X1_TC_L1D3L2D4),
.number_in_stubpair6in(SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4_number),
.read_add_stubpair6in(SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4_read_add),
.stubpair6in(SP_L1D3PHI3X1_L2D4PHI4X1_TC_L1D3L2D4),
.number_in_stubpair7in(SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4_number),
.read_add_stubpair7in(SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4_read_add),
.stubpair7in(SP_L1D3PHI1X2_L2D4PHI1X1_TC_L1D3L2D4),
.number_in_stubpair8in(SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4_number),
.read_add_stubpair8in(SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4_read_add),
.stubpair8in(SP_L1D3PHI1X2_L2D4PHI2X1_TC_L1D3L2D4),
.number_in_stubpair9in(SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4_number),
.read_add_stubpair9in(SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4_read_add),
.stubpair9in(SP_L1D3PHI2X2_L2D4PHI2X1_TC_L1D3L2D4),
.number_in_stubpair10in(SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4_number),
.read_add_stubpair10in(SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4_read_add),
.stubpair10in(SP_L1D3PHI2X2_L2D4PHI3X1_TC_L1D3L2D4),
.number_in_stubpair11in(SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4_number),
.read_add_stubpair11in(SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4_read_add),
.stubpair11in(SP_L1D3PHI3X2_L2D4PHI3X1_TC_L1D3L2D4),
.number_in_stubpair12in(SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4_number),
.read_add_stubpair12in(SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4_read_add),
.stubpair12in(SP_L1D3PHI3X2_L2D4PHI4X1_TC_L1D3L2D4),
.number_in_stubpair13in(SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4_number),
.read_add_stubpair13in(SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4_read_add),
.stubpair13in(SP_L1D3PHI1X2_L2D4PHI1X2_TC_L1D3L2D4),
.number_in_stubpair14in(SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4_number),
.read_add_stubpair14in(SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4_read_add),
.stubpair14in(SP_L1D3PHI1X2_L2D4PHI2X2_TC_L1D3L2D4),
.number_in_stubpair15in(SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4_number),
.read_add_stubpair15in(SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4_read_add),
.stubpair15in(SP_L1D3PHI2X2_L2D4PHI2X2_TC_L1D3L2D4),
.number_in_stubpair16in(SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4_number),
.read_add_stubpair16in(SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4_read_add),
.stubpair16in(SP_L1D3PHI2X2_L2D4PHI3X2_TC_L1D3L2D4),
.number_in_stubpair17in(SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4_number),
.read_add_stubpair17in(SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4_read_add),
.stubpair17in(SP_L1D3PHI3X2_L2D4PHI3X2_TC_L1D3L2D4),
.number_in_stubpair18in(SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4_number),
.read_add_stubpair18in(SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4_read_add),
.stubpair18in(SP_L1D3PHI3X2_L2D4PHI4X2_TC_L1D3L2D4),
.read_add_innerallstubin(AS_L1D3n2_TC_L1D3L2D4_read_add),
.innerallstubin(AS_L1D3n2_TC_L1D3L2D4),
.read_add_outerallstubin(AS_L2D4n1_TC_L1D3L2D4_read_add),
.outerallstubin(AS_L2D4n1_TC_L1D3L2D4),
.projoutToPlus_L3(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3),
.projoutToPlus_L4(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4),
.projoutToMinus_L3(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3),
.projoutToMinus_L4(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4),
.projout_L3D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4),
.projout_L4D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4),
.trackpar(TC_L1D3L2D4_TPAR_L1D3L2D4),
.valid_projoutToPlus_L3(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L3_wr_en),
.valid_projoutToPlus_L4(TC_L1D3L2D4_TPROJ_ToPlus_L1D3L2D4_L4_wr_en),
.valid_projoutToMinus_L3(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L3_wr_en),
.valid_projoutToMinus_L4(TC_L1D3L2D4_TPROJ_ToMinus_L1D3L2D4_L4_wr_en),
.valid_projout_L3D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L3D4_wr_en),
.valid_projout_L4D4(TC_L1D3L2D4_TPROJ_L1D3L2D4_L4D4_wr_en),
.valid_trackpar(TC_L1D3L2D4_TPAR_L1D3L2D4_wr_en),
.done_proj(TC_L1D3L2D4_proj_start),
.start(SP_L1D3PHI1X1_L2D4PHI1X1_start),
.done(TC_L1D3L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L1D3L2D3.dat"),.R1MEAN(`TC_L1L2_krA),.R2MEAN(`TC_L1L2_krB),.TC_index(4'b0010),.IsInner1(1'b1),.IsInner2(1'b1)) TC_L1D4L2D4(
.number_in_stubpair1in(SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4_number),
.read_add_stubpair1in(SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4_read_add),
.stubpair1in(SP_L1D4PHI1X1_L2D4PHI1X2_TC_L1D4L2D4),
.number_in_stubpair2in(SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4_number),
.read_add_stubpair2in(SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4_read_add),
.stubpair2in(SP_L1D4PHI1X1_L2D4PHI2X2_TC_L1D4L2D4),
.number_in_stubpair3in(SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4_number),
.read_add_stubpair3in(SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4_read_add),
.stubpair3in(SP_L1D4PHI2X1_L2D4PHI2X2_TC_L1D4L2D4),
.number_in_stubpair4in(SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4_number),
.read_add_stubpair4in(SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4_read_add),
.stubpair4in(SP_L1D4PHI2X1_L2D4PHI3X2_TC_L1D4L2D4),
.number_in_stubpair5in(SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4_number),
.read_add_stubpair5in(SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4_read_add),
.stubpair5in(SP_L1D4PHI3X1_L2D4PHI3X2_TC_L1D4L2D4),
.number_in_stubpair6in(SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4_number),
.read_add_stubpair6in(SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4_read_add),
.stubpair6in(SP_L1D4PHI3X1_L2D4PHI4X2_TC_L1D4L2D4),
.read_add_outerallstubin(AS_L2D4n2_TC_L1D4L2D4_read_add),
.outerallstubin(AS_L2D4n2_TC_L1D4L2D4),
.read_add_innerallstubin(AS_L1D4n1_TC_L1D4L2D4_read_add),
.innerallstubin(AS_L1D4n1_TC_L1D4L2D4),
.projoutToPlus_L3(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3),
.projoutToMinus_L3(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3),
.projout_L3D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4),
.trackpar(TC_L1D4L2D4_TPAR_L1D4L2D4),
.valid_projoutToPlus_L3(TC_L1D4L2D4_TPROJ_ToPlus_L1D4L2D4_L3_wr_en),
.valid_projoutToMinus_L3(TC_L1D4L2D4_TPROJ_ToMinus_L1D4L2D4_L3_wr_en),
.valid_projout_L3D4(TC_L1D4L2D4_TPROJ_L1D4L2D4_L3D4_wr_en),
.valid_trackpar(TC_L1D4L2D4_TPAR_L1D4L2D4_wr_en),
.done_proj(TC_L1D4L2D4_proj_start),
.start(SP_L1D4PHI1X1_L2D4PHI1X2_start),
.done(TC_L1D4L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L3D3L4D3.dat"),.R1MEAN(`TC_L3L4_krA),.R2MEAN(`TC_L3L4_krB),.TC_index(4'b0011),.IsInner1(1'b1),.IsInner2(1'b0)) TC_L3D3L4D3(
.number_in_stubpair1in(SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3_number),
.read_add_stubpair1in(SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3_read_add),
.stubpair1in(SP_L3D3PHI1X1_L4D3PHI1X1_TC_L3D3L4D3),
.number_in_stubpair2in(SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3_number),
.read_add_stubpair2in(SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3_read_add),
.stubpair2in(SP_L3D3PHI1X1_L4D3PHI2X1_TC_L3D3L4D3),
.number_in_stubpair3in(SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3_number),
.read_add_stubpair3in(SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3_read_add),
.stubpair3in(SP_L3D3PHI2X1_L4D3PHI2X1_TC_L3D3L4D3),
.number_in_stubpair4in(SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3_number),
.read_add_stubpair4in(SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3_read_add),
.stubpair4in(SP_L3D3PHI2X1_L4D3PHI3X1_TC_L3D3L4D3),
.number_in_stubpair5in(SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3_number),
.read_add_stubpair5in(SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3_read_add),
.stubpair5in(SP_L3D3PHI3X1_L4D3PHI3X1_TC_L3D3L4D3),
.number_in_stubpair6in(SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3_number),
.read_add_stubpair6in(SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3_read_add),
.stubpair6in(SP_L3D3PHI3X1_L4D3PHI4X1_TC_L3D3L4D3),
.number_in_stubpair7in(SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3_number),
.read_add_stubpair7in(SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3_read_add),
.stubpair7in(SP_L3D3PHI1X1_L4D3PHI1X2_TC_L3D3L4D3),
.number_in_stubpair8in(SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3_number),
.read_add_stubpair8in(SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3_read_add),
.stubpair8in(SP_L3D3PHI1X1_L4D3PHI2X2_TC_L3D3L4D3),
.number_in_stubpair9in(SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3_number),
.read_add_stubpair9in(SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3_read_add),
.stubpair9in(SP_L3D3PHI2X1_L4D3PHI2X2_TC_L3D3L4D3),
.number_in_stubpair10in(SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3_number),
.read_add_stubpair10in(SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3_read_add),
.stubpair10in(SP_L3D3PHI2X1_L4D3PHI3X2_TC_L3D3L4D3),
.number_in_stubpair11in(SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3_number),
.read_add_stubpair11in(SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3_read_add),
.stubpair11in(SP_L3D3PHI3X1_L4D3PHI3X2_TC_L3D3L4D3),
.number_in_stubpair12in(SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3_number),
.read_add_stubpair12in(SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3_read_add),
.stubpair12in(SP_L3D3PHI3X1_L4D3PHI4X2_TC_L3D3L4D3),
.number_in_stubpair13in(SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3_number),
.read_add_stubpair13in(SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3_read_add),
.stubpair13in(SP_L3D3PHI1X2_L4D3PHI1X2_TC_L3D3L4D3),
.number_in_stubpair14in(SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3_number),
.read_add_stubpair14in(SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3_read_add),
.stubpair14in(SP_L3D3PHI1X2_L4D3PHI2X2_TC_L3D3L4D3),
.number_in_stubpair15in(SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3_number),
.read_add_stubpair15in(SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3_read_add),
.stubpair15in(SP_L3D3PHI2X2_L4D3PHI2X2_TC_L3D3L4D3),
.number_in_stubpair16in(SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3_number),
.read_add_stubpair16in(SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3_read_add),
.stubpair16in(SP_L3D3PHI2X2_L4D3PHI3X2_TC_L3D3L4D3),
.number_in_stubpair17in(SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3_number),
.read_add_stubpair17in(SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3_read_add),
.stubpair17in(SP_L3D3PHI3X2_L4D3PHI3X2_TC_L3D3L4D3),
.number_in_stubpair18in(SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3_number),
.read_add_stubpair18in(SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3_read_add),
.stubpair18in(SP_L3D3PHI3X2_L4D3PHI4X2_TC_L3D3L4D3),
.read_add_outerallstubin(AS_L4D3n1_TC_L3D3L4D3_read_add),
.outerallstubin(AS_L4D3n1_TC_L3D3L4D3),
.read_add_innerallstubin(AS_L3D3n1_TC_L3D3L4D3_read_add),
.innerallstubin(AS_L3D3n1_TC_L3D3L4D3),
.projoutToPlus_L2(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2),
.projoutToPlus_L5(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5),
.projoutToPlus_L1(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1),
.projoutToPlus_L6(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6),
.projoutToMinus_L2(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2),
.projoutToMinus_L5(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5),
.projoutToMinus_L1(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1),
.projoutToMinus_L6(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6),
.projout_L1D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3),
.projout_L2D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3),
.projout_L5D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3),
.projout_L6D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3),
.projout_L5D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4),
.projout_L6D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4),
.trackpar(TC_L3D3L4D3_TPAR_L3D3L4D3),
.valid_projoutToPlus_L2(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L2_wr_en),
.valid_projoutToPlus_L5(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L5_wr_en),
.valid_projoutToPlus_L1(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L1_wr_en),
.valid_projoutToPlus_L6(TC_L3D3L4D3_TPROJ_ToPlus_L3D3L4D3_L6_wr_en),
.valid_projoutToMinus_L2(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L2_wr_en),
.valid_projoutToMinus_L5(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L5_wr_en),
.valid_projoutToMinus_L1(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L1_wr_en),
.valid_projoutToMinus_L6(TC_L3D3L4D3_TPROJ_ToMinus_L3D3L4D3_L6_wr_en),
.valid_projout_L1D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L1D3_wr_en),
.valid_projout_L2D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L2D3_wr_en),
.valid_projout_L5D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D3_wr_en),
.valid_projout_L6D3(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D3_wr_en),
.valid_projout_L5D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L5D4_wr_en),
.valid_projout_L6D4(TC_L3D3L4D3_TPROJ_L3D3L4D3_L6D4_wr_en),
.valid_trackpar(TC_L3D3L4D3_TPAR_L3D3L4D3_wr_en),
.done_proj(TC_L3D3L4D3_proj_start),
.start(SP_L3D3PHI1X1_L4D3PHI1X1_start),
.done(TC_L3D3L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L3D3L4D3.dat"),.R1MEAN(`TC_L3L4_krA),.R2MEAN(`TC_L3L4_krB),.TC_index(4'b0100),.IsInner1(1'b1),.IsInner2(1'b0)) TC_L3D3L4D4(
.number_in_stubpair1in(SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4_number),
.read_add_stubpair1in(SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4_read_add),
.stubpair1in(SP_L3D3PHI1X2_L4D4PHI1X1_TC_L3D3L4D4),
.number_in_stubpair2in(SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4_number),
.read_add_stubpair2in(SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4_read_add),
.stubpair2in(SP_L3D3PHI1X2_L4D4PHI2X1_TC_L3D3L4D4),
.number_in_stubpair3in(SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4_number),
.read_add_stubpair3in(SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4_read_add),
.stubpair3in(SP_L3D3PHI2X2_L4D4PHI2X1_TC_L3D3L4D4),
.number_in_stubpair4in(SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4_number),
.read_add_stubpair4in(SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4_read_add),
.stubpair4in(SP_L3D3PHI2X2_L4D4PHI3X1_TC_L3D3L4D4),
.number_in_stubpair5in(SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4_number),
.read_add_stubpair5in(SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4_read_add),
.stubpair5in(SP_L3D3PHI3X2_L4D4PHI3X1_TC_L3D3L4D4),
.number_in_stubpair6in(SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4_number),
.read_add_stubpair6in(SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4_read_add),
.stubpair6in(SP_L3D3PHI3X2_L4D4PHI4X1_TC_L3D3L4D4),
.read_add_innerallstubin(AS_L3D3n2_TC_L3D3L4D4_read_add),
.innerallstubin(AS_L3D3n2_TC_L3D3L4D4),
.read_add_outerallstubin(AS_L4D4n1_TC_L3D3L4D4_read_add),
.outerallstubin(AS_L4D4n1_TC_L3D3L4D4),
.projoutToPlus_L2(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2),
.projoutToPlus_L5(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5),
.projoutToPlus_L1(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1),
.projoutToPlus_L6(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6),
.projoutToMinus_L2(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2),
.projoutToMinus_L5(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5),
.projoutToMinus_L1(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1),
.projoutToMinus_L6(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6),
.projout_L1D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3),
.projout_L2D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3),
.projout_L5D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4),
.projout_L6D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4),
.trackpar(TC_L3D3L4D4_TPAR_L3D3L4D4),
.valid_projoutToPlus_L2(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L2_wr_en),
.valid_projoutToPlus_L5(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L5_wr_en),
.valid_projoutToPlus_L1(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L1_wr_en),
.valid_projoutToPlus_L6(TC_L3D3L4D4_TPROJ_ToPlus_L3D3L4D4_L6_wr_en),
.valid_projoutToMinus_L2(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L2_wr_en),
.valid_projoutToMinus_L5(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L5_wr_en),
.valid_projoutToMinus_L1(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L1_wr_en),
.valid_projoutToMinus_L6(TC_L3D3L4D4_TPROJ_ToMinus_L3D3L4D4_L6_wr_en),
.valid_projout_L1D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L1D3_wr_en),
.valid_projout_L2D3(TC_L3D3L4D4_TPROJ_L3D3L4D4_L2D3_wr_en),
.valid_projout_L5D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L5D4_wr_en),
.valid_projout_L6D4(TC_L3D3L4D4_TPROJ_L3D3L4D4_L6D4_wr_en),
.valid_trackpar(TC_L3D3L4D4_TPAR_L3D3L4D4_wr_en),
.done_proj(TC_L3D3L4D4_proj_start),
.start(SP_L3D3PHI1X2_L4D4PHI1X1_start),
.done(TC_L3D3L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L3D3L4D3.dat"),.R1MEAN(`TC_L3L4_krA),.R2MEAN(`TC_L3L4_krB),.TC_index(4'b0101),.IsInner1(1'b1),.IsInner2(1'b0)) TC_L3D4L4D4(
.number_in_stubpair1in(SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4_number),
.read_add_stubpair1in(SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4_read_add),
.stubpair1in(SP_L3D4PHI1X1_L4D4PHI1X1_TC_L3D4L4D4),
.number_in_stubpair2in(SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4_number),
.read_add_stubpair2in(SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4_read_add),
.stubpair2in(SP_L3D4PHI1X1_L4D4PHI2X1_TC_L3D4L4D4),
.number_in_stubpair3in(SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4_number),
.read_add_stubpair3in(SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4_read_add),
.stubpair3in(SP_L3D4PHI2X1_L4D4PHI2X1_TC_L3D4L4D4),
.number_in_stubpair4in(SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4_number),
.read_add_stubpair4in(SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4_read_add),
.stubpair4in(SP_L3D4PHI2X1_L4D4PHI3X1_TC_L3D4L4D4),
.number_in_stubpair5in(SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4_number),
.read_add_stubpair5in(SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4_read_add),
.stubpair5in(SP_L3D4PHI3X1_L4D4PHI3X1_TC_L3D4L4D4),
.number_in_stubpair6in(SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4_number),
.read_add_stubpair6in(SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4_read_add),
.stubpair6in(SP_L3D4PHI3X1_L4D4PHI4X1_TC_L3D4L4D4),
.number_in_stubpair7in(SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4_number),
.read_add_stubpair7in(SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4_read_add),
.stubpair7in(SP_L3D4PHI1X1_L4D4PHI1X2_TC_L3D4L4D4),
.number_in_stubpair8in(SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4_number),
.read_add_stubpair8in(SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4_read_add),
.stubpair8in(SP_L3D4PHI1X1_L4D4PHI2X2_TC_L3D4L4D4),
.number_in_stubpair9in(SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4_number),
.read_add_stubpair9in(SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4_read_add),
.stubpair9in(SP_L3D4PHI2X1_L4D4PHI2X2_TC_L3D4L4D4),
.number_in_stubpair10in(SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4_number),
.read_add_stubpair10in(SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4_read_add),
.stubpair10in(SP_L3D4PHI2X1_L4D4PHI3X2_TC_L3D4L4D4),
.number_in_stubpair11in(SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4_number),
.read_add_stubpair11in(SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4_read_add),
.stubpair11in(SP_L3D4PHI3X1_L4D4PHI3X2_TC_L3D4L4D4),
.number_in_stubpair12in(SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4_number),
.read_add_stubpair12in(SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4_read_add),
.stubpair12in(SP_L3D4PHI3X1_L4D4PHI4X2_TC_L3D4L4D4),
.number_in_stubpair13in(SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4_number),
.read_add_stubpair13in(SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4_read_add),
.stubpair13in(SP_L3D4PHI1X2_L4D4PHI1X2_TC_L3D4L4D4),
.number_in_stubpair14in(SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4_number),
.read_add_stubpair14in(SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4_read_add),
.stubpair14in(SP_L3D4PHI1X2_L4D4PHI2X2_TC_L3D4L4D4),
.number_in_stubpair15in(SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4_number),
.read_add_stubpair15in(SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4_read_add),
.stubpair15in(SP_L3D4PHI2X2_L4D4PHI2X2_TC_L3D4L4D4),
.number_in_stubpair16in(SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4_number),
.read_add_stubpair16in(SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4_read_add),
.stubpair16in(SP_L3D4PHI2X2_L4D4PHI3X2_TC_L3D4L4D4),
.number_in_stubpair17in(SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4_number),
.read_add_stubpair17in(SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4_read_add),
.stubpair17in(SP_L3D4PHI3X2_L4D4PHI3X2_TC_L3D4L4D4),
.number_in_stubpair18in(SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4_number),
.read_add_stubpair18in(SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4_read_add),
.stubpair18in(SP_L3D4PHI3X2_L4D4PHI4X2_TC_L3D4L4D4),
.read_add_outerallstubin(AS_L4D4n2_TC_L3D4L4D4_read_add),
.outerallstubin(AS_L4D4n2_TC_L3D4L4D4),
.read_add_innerallstubin(AS_L3D4n1_TC_L3D4L4D4_read_add),
.innerallstubin(AS_L3D4n1_TC_L3D4L4D4),
.projoutToPlus_L2(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2),
.projoutToPlus_L5(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5),
.projoutToPlus_L1(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1),
.projoutToPlus_L6(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6),
.projoutToMinus_L2(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2),
.projoutToMinus_L5(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5),
.projoutToMinus_L1(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1),
.projoutToMinus_L6(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6),
.projout_L1D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3),
.projout_L2D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3),
.projout_L2D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4),
.projout_L5D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4),
.projout_L6D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4),
.trackpar(TC_L3D4L4D4_TPAR_L3D4L4D4),
.valid_projoutToPlus_L2(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L2_wr_en),
.valid_projoutToPlus_L5(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L5_wr_en),
.valid_projoutToPlus_L1(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L1_wr_en),
.valid_projoutToPlus_L6(TC_L3D4L4D4_TPROJ_ToPlus_L3D4L4D4_L6_wr_en),
.valid_projoutToMinus_L2(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L2_wr_en),
.valid_projoutToMinus_L5(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L5_wr_en),
.valid_projoutToMinus_L1(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L1_wr_en),
.valid_projoutToMinus_L6(TC_L3D4L4D4_TPROJ_ToMinus_L3D4L4D4_L6_wr_en),
.valid_projout_L1D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L1D3_wr_en),
.valid_projout_L2D3(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D3_wr_en),
.valid_projout_L2D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L2D4_wr_en),
.valid_projout_L5D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L5D4_wr_en),
.valid_projout_L6D4(TC_L3D4L4D4_TPROJ_L3D4L4D4_L6D4_wr_en),
.valid_trackpar(TC_L3D4L4D4_TPAR_L3D4L4D4_wr_en),
.done_proj(TC_L3D4L4D4_proj_start),
.start(SP_L3D4PHI1X1_L4D4PHI1X1_start),
.done(TC_L3D4L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L5D3L6D3.dat"),.R1MEAN(`TC_L5L6_krA),.R2MEAN(`TC_L5L6_krB),.TC_index(4'b0011),.IsInner1(1'b0),.IsInner2(1'b0)) TC_L5D3L6D3(
.number_in_stubpair1in(SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3_number),
.read_add_stubpair1in(SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3_read_add),
.stubpair1in(SP_L5D3PHI1X1_L6D3PHI1X1_TC_L5D3L6D3),
.number_in_stubpair2in(SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3_number),
.read_add_stubpair2in(SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3_read_add),
.stubpair2in(SP_L5D3PHI1X1_L6D3PHI2X1_TC_L5D3L6D3),
.number_in_stubpair3in(SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3_number),
.read_add_stubpair3in(SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3_read_add),
.stubpair3in(SP_L5D3PHI2X1_L6D3PHI2X1_TC_L5D3L6D3),
.number_in_stubpair4in(SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3_number),
.read_add_stubpair4in(SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3_read_add),
.stubpair4in(SP_L5D3PHI2X1_L6D3PHI3X1_TC_L5D3L6D3),
.number_in_stubpair5in(SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3_number),
.read_add_stubpair5in(SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3_read_add),
.stubpair5in(SP_L5D3PHI3X1_L6D3PHI3X1_TC_L5D3L6D3),
.number_in_stubpair6in(SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3_number),
.read_add_stubpair6in(SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3_read_add),
.stubpair6in(SP_L5D3PHI3X1_L6D3PHI4X1_TC_L5D3L6D3),
.number_in_stubpair7in(SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3_number),
.read_add_stubpair7in(SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3_read_add),
.stubpair7in(SP_L5D3PHI1X1_L6D3PHI1X2_TC_L5D3L6D3),
.number_in_stubpair8in(SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3_number),
.read_add_stubpair8in(SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3_read_add),
.stubpair8in(SP_L5D3PHI1X1_L6D3PHI2X2_TC_L5D3L6D3),
.number_in_stubpair9in(SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3_number),
.read_add_stubpair9in(SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3_read_add),
.stubpair9in(SP_L5D3PHI2X1_L6D3PHI2X2_TC_L5D3L6D3),
.number_in_stubpair10in(SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3_number),
.read_add_stubpair10in(SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3_read_add),
.stubpair10in(SP_L5D3PHI2X1_L6D3PHI3X2_TC_L5D3L6D3),
.number_in_stubpair11in(SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3_number),
.read_add_stubpair11in(SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3_read_add),
.stubpair11in(SP_L5D3PHI3X1_L6D3PHI3X2_TC_L5D3L6D3),
.number_in_stubpair12in(SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3_number),
.read_add_stubpair12in(SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3_read_add),
.stubpair12in(SP_L5D3PHI3X1_L6D3PHI4X2_TC_L5D3L6D3),
.number_in_stubpair13in(SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3_number),
.read_add_stubpair13in(SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3_read_add),
.stubpair13in(SP_L5D3PHI1X2_L6D3PHI1X2_TC_L5D3L6D3),
.number_in_stubpair14in(SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3_number),
.read_add_stubpair14in(SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3_read_add),
.stubpair14in(SP_L5D3PHI1X2_L6D3PHI2X2_TC_L5D3L6D3),
.number_in_stubpair15in(SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3_number),
.read_add_stubpair15in(SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3_read_add),
.stubpair15in(SP_L5D3PHI2X2_L6D3PHI2X2_TC_L5D3L6D3),
.number_in_stubpair16in(SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3_number),
.read_add_stubpair16in(SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3_read_add),
.stubpair16in(SP_L5D3PHI2X2_L6D3PHI3X2_TC_L5D3L6D3),
.number_in_stubpair17in(SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3_number),
.read_add_stubpair17in(SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3_read_add),
.stubpair17in(SP_L5D3PHI3X2_L6D3PHI3X2_TC_L5D3L6D3),
.number_in_stubpair18in(SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3_number),
.read_add_stubpair18in(SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3_read_add),
.stubpair18in(SP_L5D3PHI3X2_L6D3PHI4X2_TC_L5D3L6D3),
.read_add_outerallstubin(AS_L6D3n1_TC_L5D3L6D3_read_add),
.outerallstubin(AS_L6D3n1_TC_L5D3L6D3),
.read_add_innerallstubin(AS_L5D3n1_TC_L5D3L6D3_read_add),
.innerallstubin(AS_L5D3n1_TC_L5D3L6D3),
.projoutToPlus_L3(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3),
.projoutToPlus_L4(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4),
.projoutToPlus_L2(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2),
.projoutToPlus_L1(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1),
.projoutToMinus_L3(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3),
.projoutToMinus_L4(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4),
.projoutToMinus_L2(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2),
.projoutToMinus_L1(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1),
.projout_L1D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3),
.projout_L2D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3),
.projout_L3D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3),
.projout_L4D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3),
.trackpar(TC_L5D3L6D3_TPAR_L5D3L6D3),
.valid_projoutToPlus_L3(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L3_wr_en),
.valid_projoutToPlus_L4(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L4_wr_en),
.valid_projoutToPlus_L2(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L2_wr_en),
.valid_projoutToPlus_L1(TC_L5D3L6D3_TPROJ_ToPlus_L5D3L6D3_L1_wr_en),
.valid_projoutToMinus_L3(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L3_wr_en),
.valid_projoutToMinus_L4(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L4_wr_en),
.valid_projoutToMinus_L2(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L2_wr_en),
.valid_projoutToMinus_L1(TC_L5D3L6D3_TPROJ_ToMinus_L5D3L6D3_L1_wr_en),
.valid_projout_L1D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L1D3_wr_en),
.valid_projout_L2D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L2D3_wr_en),
.valid_projout_L3D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L3D3_wr_en),
.valid_projout_L4D3(TC_L5D3L6D3_TPROJ_L5D3L6D3_L4D3_wr_en),
.valid_trackpar(TC_L5D3L6D3_TPAR_L5D3L6D3_wr_en),
.done_proj(TC_L5D3L6D3_proj_start),
.start(SP_L5D3PHI1X1_L6D3PHI1X1_start),
.done(TC_L5D3L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L5D3L6D3.dat"),.R1MEAN(`TC_L5L6_krA),.R2MEAN(`TC_L5L6_krB),.TC_index(4'b0100),.IsInner1(1'b0),.IsInner2(1'b0)) TC_L5D3L6D4(
.number_in_stubpair1in(SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4_number),
.read_add_stubpair1in(SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4_read_add),
.stubpair1in(SP_L5D3PHI1X2_L6D4PHI1X1_TC_L5D3L6D4),
.number_in_stubpair2in(SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4_number),
.read_add_stubpair2in(SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4_read_add),
.stubpair2in(SP_L5D3PHI1X2_L6D4PHI2X1_TC_L5D3L6D4),
.number_in_stubpair3in(SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4_number),
.read_add_stubpair3in(SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4_read_add),
.stubpair3in(SP_L5D3PHI2X2_L6D4PHI2X1_TC_L5D3L6D4),
.number_in_stubpair4in(SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4_number),
.read_add_stubpair4in(SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4_read_add),
.stubpair4in(SP_L5D3PHI2X2_L6D4PHI3X1_TC_L5D3L6D4),
.number_in_stubpair5in(SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4_number),
.read_add_stubpair5in(SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4_read_add),
.stubpair5in(SP_L5D3PHI3X2_L6D4PHI3X1_TC_L5D3L6D4),
.number_in_stubpair6in(SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4_number),
.read_add_stubpair6in(SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4_read_add),
.stubpair6in(SP_L5D3PHI3X2_L6D4PHI4X1_TC_L5D3L6D4),
.read_add_innerallstubin(AS_L5D3n2_TC_L5D3L6D4_read_add),
.innerallstubin(AS_L5D3n2_TC_L5D3L6D4),
.read_add_outerallstubin(AS_L6D4n1_TC_L5D3L6D4_read_add),
.outerallstubin(AS_L6D4n1_TC_L5D3L6D4),
.projoutToPlus_L3(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3),
.projoutToPlus_L4(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4),
.projoutToPlus_L2(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2),
.projoutToPlus_L1(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1),
.projoutToMinus_L3(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3),
.projoutToMinus_L4(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4),
.projoutToMinus_L2(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2),
.projoutToMinus_L1(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1),
.projout_L1D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3),
.projout_L2D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3),
.projout_L3D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3),
.projout_L4D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3),
.trackpar(TC_L5D3L6D4_TPAR_L5D3L6D4),
.valid_projoutToPlus_L3(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L3_wr_en),
.valid_projoutToPlus_L4(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L4_wr_en),
.valid_projoutToPlus_L2(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L2_wr_en),
.valid_projoutToPlus_L1(TC_L5D3L6D4_TPROJ_ToPlus_L5D3L6D4_L1_wr_en),
.valid_projoutToMinus_L3(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L3_wr_en),
.valid_projoutToMinus_L4(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L4_wr_en),
.valid_projoutToMinus_L2(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L2_wr_en),
.valid_projoutToMinus_L1(TC_L5D3L6D4_TPROJ_ToMinus_L5D3L6D4_L1_wr_en),
.valid_projout_L1D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L1D3_wr_en),
.valid_projout_L2D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L2D3_wr_en),
.valid_projout_L3D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L3D3_wr_en),
.valid_projout_L4D3(TC_L5D3L6D4_TPROJ_L5D3L6D4_L4D3_wr_en),
.valid_trackpar(TC_L5D3L6D4_TPAR_L5D3L6D4_wr_en),
.done_proj(TC_L5D3L6D4_proj_start),
.start(SP_L5D3PHI1X2_L6D4PHI1X1_start),
.done(TC_L5D3L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

TrackletCalculator #(.BARREL(1'b1),.InvR_FILE("InvRTable_TC_L5D3L6D3.dat"),.R1MEAN(`TC_L5L6_krA),.R2MEAN(`TC_L5L6_krB),.TC_index(4'b0101),.IsInner1(1'b0),.IsInner2(1'b0)) TC_L5D4L6D4(
.number_in_stubpair1in(SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4_number),
.read_add_stubpair1in(SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4_read_add),
.stubpair1in(SP_L5D4PHI1X1_L6D4PHI1X1_TC_L5D4L6D4),
.number_in_stubpair2in(SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4_number),
.read_add_stubpair2in(SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4_read_add),
.stubpair2in(SP_L5D4PHI1X1_L6D4PHI2X1_TC_L5D4L6D4),
.number_in_stubpair3in(SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4_number),
.read_add_stubpair3in(SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4_read_add),
.stubpair3in(SP_L5D4PHI2X1_L6D4PHI2X1_TC_L5D4L6D4),
.number_in_stubpair4in(SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4_number),
.read_add_stubpair4in(SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4_read_add),
.stubpair4in(SP_L5D4PHI2X1_L6D4PHI3X1_TC_L5D4L6D4),
.number_in_stubpair5in(SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4_number),
.read_add_stubpair5in(SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4_read_add),
.stubpair5in(SP_L5D4PHI3X1_L6D4PHI3X1_TC_L5D4L6D4),
.number_in_stubpair6in(SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4_number),
.read_add_stubpair6in(SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4_read_add),
.stubpair6in(SP_L5D4PHI3X1_L6D4PHI4X1_TC_L5D4L6D4),
.number_in_stubpair7in(SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4_number),
.read_add_stubpair7in(SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4_read_add),
.stubpair7in(SP_L5D4PHI1X1_L6D4PHI1X2_TC_L5D4L6D4),
.number_in_stubpair8in(SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4_number),
.read_add_stubpair8in(SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4_read_add),
.stubpair8in(SP_L5D4PHI1X1_L6D4PHI2X2_TC_L5D4L6D4),
.number_in_stubpair9in(SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4_number),
.read_add_stubpair9in(SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4_read_add),
.stubpair9in(SP_L5D4PHI2X1_L6D4PHI2X2_TC_L5D4L6D4),
.number_in_stubpair10in(SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4_number),
.read_add_stubpair10in(SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4_read_add),
.stubpair10in(SP_L5D4PHI2X1_L6D4PHI3X2_TC_L5D4L6D4),
.number_in_stubpair11in(SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4_number),
.read_add_stubpair11in(SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4_read_add),
.stubpair11in(SP_L5D4PHI3X1_L6D4PHI3X2_TC_L5D4L6D4),
.number_in_stubpair12in(SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4_number),
.read_add_stubpair12in(SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4_read_add),
.stubpair12in(SP_L5D4PHI3X1_L6D4PHI4X2_TC_L5D4L6D4),
.number_in_stubpair13in(SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4_number),
.read_add_stubpair13in(SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4_read_add),
.stubpair13in(SP_L5D4PHI1X2_L6D4PHI1X2_TC_L5D4L6D4),
.number_in_stubpair14in(SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4_number),
.read_add_stubpair14in(SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4_read_add),
.stubpair14in(SP_L5D4PHI1X2_L6D4PHI2X2_TC_L5D4L6D4),
.number_in_stubpair15in(SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4_number),
.read_add_stubpair15in(SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4_read_add),
.stubpair15in(SP_L5D4PHI2X2_L6D4PHI2X2_TC_L5D4L6D4),
.number_in_stubpair16in(SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4_number),
.read_add_stubpair16in(SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4_read_add),
.stubpair16in(SP_L5D4PHI2X2_L6D4PHI3X2_TC_L5D4L6D4),
.number_in_stubpair17in(SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4_number),
.read_add_stubpair17in(SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4_read_add),
.stubpair17in(SP_L5D4PHI3X2_L6D4PHI3X2_TC_L5D4L6D4),
.number_in_stubpair18in(SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4_number),
.read_add_stubpair18in(SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4_read_add),
.stubpair18in(SP_L5D4PHI3X2_L6D4PHI4X2_TC_L5D4L6D4),
.read_add_outerallstubin(AS_L6D4n2_TC_L5D4L6D4_read_add),
.outerallstubin(AS_L6D4n2_TC_L5D4L6D4),
.read_add_innerallstubin(AS_L5D4n1_TC_L5D4L6D4_read_add),
.innerallstubin(AS_L5D4n1_TC_L5D4L6D4),
.projoutToPlus_L3(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3),
.projoutToPlus_L4(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4),
.projoutToPlus_L2(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2),
.projoutToPlus_L1(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1),
.projoutToMinus_L3(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3),
.projoutToMinus_L4(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4),
.projoutToMinus_L2(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2),
.projoutToMinus_L1(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1),
.projout_L1D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3),
.projout_L2D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3),
.projout_L3D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3),
.projout_L4D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3),
.projout_L3D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4),
.projout_L4D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4),
.trackpar(TC_L5D4L6D4_TPAR_L5D4L6D4),
.valid_projoutToPlus_L3(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L3_wr_en),
.valid_projoutToPlus_L4(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L4_wr_en),
.valid_projoutToPlus_L2(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L2_wr_en),
.valid_projoutToPlus_L1(TC_L5D4L6D4_TPROJ_ToPlus_L5D4L6D4_L1_wr_en),
.valid_projoutToMinus_L3(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L3_wr_en),
.valid_projoutToMinus_L4(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L4_wr_en),
.valid_projoutToMinus_L2(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L2_wr_en),
.valid_projoutToMinus_L1(TC_L5D4L6D4_TPROJ_ToMinus_L5D4L6D4_L1_wr_en),
.valid_projout_L1D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L1D3_wr_en),
.valid_projout_L2D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L2D3_wr_en),
.valid_projout_L3D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D3_wr_en),
.valid_projout_L4D3(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D3_wr_en),
.valid_projout_L3D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L3D4_wr_en),
.valid_projout_L4D4(TC_L5D4L6D4_TPROJ_L5D4L6D4_L4D4_wr_en),
.valid_trackpar(TC_L5D4L6D4_TPAR_L5D4L6D4_wr_en),
.done_proj(TC_L5D4L6D4_proj_start),
.start(SP_L5D4PHI1X1_L6D4PHI1X1_start),
.done(TC_L5D4L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L3F3F5") PT_L3F3F5_Plus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus_number),
.read_add_projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus_read_add),
.projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L3_PT_L3F3F5_Plus),
.number_in_projin_layer_2(TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus_number),
.read_add_projin_layer_2(TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus_read_add),
.projin_layer_2(TPROJ_ToPlus_L1D3L2D4_L3_PT_L3F3F5_Plus),
.number_in_projin_layer_3(TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus_number),
.read_add_projin_layer_3(TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus_read_add),
.projin_layer_3(TPROJ_ToPlus_L1D4L2D4_L3_PT_L3F3F5_Plus),
.number_in_projin_layer_4(TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus_number),
.read_add_projin_layer_4(TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus_read_add),
.projin_layer_4(TPROJ_ToPlus_L5D3L6D3_L3_PT_L3F3F5_Plus),
.number_in_projin_layer_5(TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus_number),
.read_add_projin_layer_5(TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus_read_add),
.projin_layer_5(TPROJ_ToPlus_L5D3L6D4_L3_PT_L3F3F5_Plus),
.number_in_projin_layer_6(TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus_number),
.read_add_projin_layer_6(TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus_read_add),
.projin_layer_6(TPROJ_ToPlus_L5D4L6D4_L3_PT_L3F3F5_Plus),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L3F3F5_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L3F3F5_Plus_From_DataStream),
.projout_layer_1(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L1L2),
.valid_layer_1(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L1L2_wr_en),
.projout_layer_2(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L1L2),
.valid_layer_2(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L1L2_wr_en),
.projout_layer_3(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L5L6),
.valid_layer_3(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D3_L5L6_wr_en),
.projout_layer_4(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L5L6),
.valid_layer_4(PT_L3F3F5_Plus_TPROJ_FromPlus_L3D4_L5L6_wr_en),
.valid_proj_data_stream(PT_L3F3F5_Plus_To_DataStream_en),
.proj_data_stream(PT_L3F3F5_Plus_To_DataStream),
.start(TPROJ_ToPlus_L5D4L6D4_L3_start),
.done(PT_L3F3F5_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L2L4F2") PT_L2L4F2_Plus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus_number),
.read_add_projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus_read_add),
.projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L4_PT_L2L4F2_Plus),
.number_in_projin_layer_2(TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus_number),
.read_add_projin_layer_2(TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus_read_add),
.projin_layer_2(TPROJ_ToPlus_L1D3L2D4_L4_PT_L2L4F2_Plus),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus_number),
.read_add_projin_layer_4(TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus_read_add),
.projin_layer_4(TPROJ_ToPlus_L5D3L6D3_L4_PT_L2L4F2_Plus),
.number_in_projin_layer_5(TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus_number),
.read_add_projin_layer_5(TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus_read_add),
.projin_layer_5(TPROJ_ToPlus_L5D3L6D4_L4_PT_L2L4F2_Plus),
.number_in_projin_layer_6(TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus_number),
.read_add_projin_layer_6(TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus_read_add),
.projin_layer_6(TPROJ_ToPlus_L5D4L6D4_L4_PT_L2L4F2_Plus),
.number_in_projin_layer_7(TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus_number),
.read_add_projin_layer_7(TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus_read_add),
.projin_layer_7(TPROJ_ToPlus_L3D3L4D3_L2_PT_L2L4F2_Plus),
.number_in_projin_layer_8(TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus_number),
.read_add_projin_layer_8(TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus_read_add),
.projin_layer_8(TPROJ_ToPlus_L3D3L4D4_L2_PT_L2L4F2_Plus),
.number_in_projin_layer_9(TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus_number),
.read_add_projin_layer_9(TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus_read_add),
.projin_layer_9(TPROJ_ToPlus_L3D4L4D4_L2_PT_L2L4F2_Plus),
.number_in_projin_layer_10(TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus_number),
.read_add_projin_layer_10(TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus_read_add),
.projin_layer_10(TPROJ_ToPlus_L5D3L6D3_L2_PT_L2L4F2_Plus),
.number_in_projin_layer_11(TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus_number),
.read_add_projin_layer_11(TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus_read_add),
.projin_layer_11(TPROJ_ToPlus_L5D3L6D4_L2_PT_L2L4F2_Plus),
.number_in_projin_layer_12(TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus_number),
.read_add_projin_layer_12(TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus_read_add),
.projin_layer_12(TPROJ_ToPlus_L5D4L6D4_L2_PT_L2L4F2_Plus),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L2L4F2_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L2L4F2_Plus_From_DataStream),
.projout_layer_1(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L3L4),
.valid_layer_1(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L3L4_wr_en),
.projout_layer_2(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L3L4),
.valid_layer_2(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L3L4_wr_en),
.projout_layer_3(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L1L2),
.valid_layer_3(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L1L2_wr_en),
.projout_layer_4(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L1L2),
.valid_layer_4(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L1L2_wr_en),
.projout_layer_5(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L5L6),
.valid_layer_5(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D3_L5L6_wr_en),
.projout_layer_6(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L5L6),
.valid_layer_6(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D3_L5L6_wr_en),
.projout_layer_7(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L5L6),
.valid_layer_7(PT_L2L4F2_Plus_TPROJ_FromPlus_L2D4_L5L6_wr_en),
.projout_layer_8(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L5L6),
.valid_layer_8(PT_L2L4F2_Plus_TPROJ_FromPlus_L4D4_L5L6_wr_en),
.valid_proj_data_stream(PT_L2L4F2_Plus_To_DataStream_en),
.proj_data_stream(PT_L2L4F2_Plus_To_DataStream),
.start(TPROJ_ToPlus_L5D4L6D4_L4_start),
.done(PT_L2L4F2_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("F1L5") PT_F1L5_Plus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus_number),
.read_add_projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus_read_add),
.projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L5_PT_F1L5_Plus),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus_number),
.read_add_projin_layer_4(TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus_read_add),
.projin_layer_4(TPROJ_ToPlus_L3D3L4D3_L5_PT_F1L5_Plus),
.number_in_projin_layer_5(TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus_number),
.read_add_projin_layer_5(TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus_read_add),
.projin_layer_5(TPROJ_ToPlus_L3D3L4D4_L5_PT_F1L5_Plus),
.number_in_projin_layer_6(TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus_number),
.read_add_projin_layer_6(TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus_read_add),
.projin_layer_6(TPROJ_ToPlus_L3D4L4D4_L5_PT_F1L5_Plus),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_F1L5_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_F1L5_Plus_From_DataStream),
.projout_layer_1(PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L3L4),
.valid_layer_1(PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L3L4_wr_en),
.projout_layer_2(PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L3L4),
.valid_layer_2(PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L3L4_wr_en),
.projout_layer_3(PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L1L2),
.valid_layer_3(PT_F1L5_Plus_TPROJ_FromPlus_L5D3_L1L2_wr_en),
.projout_layer_4(PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L1L2),
.valid_layer_4(PT_F1L5_Plus_TPROJ_FromPlus_L5D4_L1L2_wr_en),
.valid_proj_data_stream(PT_F1L5_Plus_To_DataStream_en),
.proj_data_stream(PT_F1L5_Plus_To_DataStream),
.start(TPROJ_ToPlus_L3D4L4D4_L5_start),
.done(PT_F1L5_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L1L6F4") PT_L1L6F4_Plus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus_number),
.read_add_projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus_read_add),
.projin_layer_1(TPROJ_ToPlus_L1D3L2D3_L6_PT_L1L6F4_Plus),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus_number),
.read_add_projin_layer_4(TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus_read_add),
.projin_layer_4(TPROJ_ToPlus_L3D3L4D3_L6_PT_L1L6F4_Plus),
.number_in_projin_layer_5(TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus_number),
.read_add_projin_layer_5(TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus_read_add),
.projin_layer_5(TPROJ_ToPlus_L3D3L4D4_L6_PT_L1L6F4_Plus),
.number_in_projin_layer_6(TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus_number),
.read_add_projin_layer_6(TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus_read_add),
.projin_layer_6(TPROJ_ToPlus_L3D4L4D4_L6_PT_L1L6F4_Plus),
.number_in_projin_layer_7(TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus_number),
.read_add_projin_layer_7(TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus_read_add),
.projin_layer_7(TPROJ_ToPlus_L3D3L4D3_L1_PT_L1L6F4_Plus),
.number_in_projin_layer_8(TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus_number),
.read_add_projin_layer_8(TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus_read_add),
.projin_layer_8(TPROJ_ToPlus_L3D3L4D4_L1_PT_L1L6F4_Plus),
.number_in_projin_layer_9(TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus_number),
.read_add_projin_layer_9(TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus_read_add),
.projin_layer_9(TPROJ_ToPlus_L3D4L4D4_L1_PT_L1L6F4_Plus),
.number_in_projin_layer_10(TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus_number),
.read_add_projin_layer_10(TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus_read_add),
.projin_layer_10(TPROJ_ToPlus_L5D3L6D3_L1_PT_L1L6F4_Plus),
.number_in_projin_layer_11(TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus_number),
.read_add_projin_layer_11(TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus_read_add),
.projin_layer_11(TPROJ_ToPlus_L5D3L6D4_L1_PT_L1L6F4_Plus),
.number_in_projin_layer_12(TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus_number),
.read_add_projin_layer_12(TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus_read_add),
.projin_layer_12(TPROJ_ToPlus_L5D4L6D4_L1_PT_L1L6F4_Plus),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L1L6F4_Plus_From_DataStream_en),
.incomming_proj_data_stream(PT_L1L6F4_Plus_From_DataStream),
.projout_layer_1(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L3L4),
.valid_layer_1(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L3L4_wr_en),
.projout_layer_2(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L3L4),
.valid_layer_2(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L3L4_wr_en),
.projout_layer_3(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L3L4),
.valid_layer_3(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L3L4_wr_en),
.projout_layer_4(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L3L4),
.valid_layer_4(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L3L4_wr_en),
.projout_layer_5(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L1L2),
.valid_layer_5(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D3_L1L2_wr_en),
.projout_layer_6(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L1L2),
.valid_layer_6(PT_L1L6F4_Plus_TPROJ_FromPlus_L6D4_L1L2_wr_en),
.projout_layer_7(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L5L6),
.valid_layer_7(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D3_L5L6_wr_en),
.projout_layer_8(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L5L6),
.valid_layer_8(PT_L1L6F4_Plus_TPROJ_FromPlus_L1D4_L5L6_wr_en),
.valid_proj_data_stream(PT_L1L6F4_Plus_To_DataStream_en),
.proj_data_stream(PT_L1L6F4_Plus_To_DataStream),
.start(TPROJ_ToPlus_L5D4L6D4_L1_start),
.done(PT_L1L6F4_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L3F3F5") PT_L3F3F5_Minus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus_number),
.read_add_projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus_read_add),
.projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L3_PT_L3F3F5_Minus),
.number_in_projin_layer_2(TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus_number),
.read_add_projin_layer_2(TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus_read_add),
.projin_layer_2(TPROJ_ToMinus_L1D3L2D4_L3_PT_L3F3F5_Minus),
.number_in_projin_layer_3(TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus_number),
.read_add_projin_layer_3(TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus_read_add),
.projin_layer_3(TPROJ_ToMinus_L1D4L2D4_L3_PT_L3F3F5_Minus),
.number_in_projin_layer_4(TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus_number),
.read_add_projin_layer_4(TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus_read_add),
.projin_layer_4(TPROJ_ToMinus_L5D3L6D3_L3_PT_L3F3F5_Minus),
.number_in_projin_layer_5(TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus_number),
.read_add_projin_layer_5(TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus_read_add),
.projin_layer_5(TPROJ_ToMinus_L5D3L6D4_L3_PT_L3F3F5_Minus),
.number_in_projin_layer_6(TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus_number),
.read_add_projin_layer_6(TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus_read_add),
.projin_layer_6(TPROJ_ToMinus_L5D4L6D4_L3_PT_L3F3F5_Minus),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L3F3F5_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L3F3F5_Minus_From_DataStream),
.projout_layer_1(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L1L2),
.valid_layer_1(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L1L2_wr_en),
.projout_layer_2(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L1L2),
.valid_layer_2(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L1L2_wr_en),
.projout_layer_3(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L5L6),
.valid_layer_3(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D3_L5L6_wr_en),
.projout_layer_4(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L5L6),
.valid_layer_4(PT_L3F3F5_Minus_TPROJ_FromMinus_L3D4_L5L6_wr_en),
.valid_proj_data_stream(PT_L3F3F5_Minus_To_DataStream_en),
.proj_data_stream(PT_L3F3F5_Minus_To_DataStream),
.start(TPROJ_ToMinus_L5D4L6D4_L3_start),
.done(PT_L3F3F5_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L2L4F2") PT_L2L4F2_Minus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus_number),
.read_add_projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus_read_add),
.projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L4_PT_L2L4F2_Minus),
.number_in_projin_layer_2(TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus_number),
.read_add_projin_layer_2(TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus_read_add),
.projin_layer_2(TPROJ_ToMinus_L1D3L2D4_L4_PT_L2L4F2_Minus),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus_number),
.read_add_projin_layer_4(TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus_read_add),
.projin_layer_4(TPROJ_ToMinus_L5D3L6D3_L4_PT_L2L4F2_Minus),
.number_in_projin_layer_5(TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus_number),
.read_add_projin_layer_5(TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus_read_add),
.projin_layer_5(TPROJ_ToMinus_L5D3L6D4_L4_PT_L2L4F2_Minus),
.number_in_projin_layer_6(TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus_number),
.read_add_projin_layer_6(TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus_read_add),
.projin_layer_6(TPROJ_ToMinus_L5D4L6D4_L4_PT_L2L4F2_Minus),
.number_in_projin_layer_7(TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus_number),
.read_add_projin_layer_7(TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus_read_add),
.projin_layer_7(TPROJ_ToMinus_L3D3L4D3_L2_PT_L2L4F2_Minus),
.number_in_projin_layer_8(TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus_number),
.read_add_projin_layer_8(TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus_read_add),
.projin_layer_8(TPROJ_ToMinus_L3D3L4D4_L2_PT_L2L4F2_Minus),
.number_in_projin_layer_9(TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus_number),
.read_add_projin_layer_9(TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus_read_add),
.projin_layer_9(TPROJ_ToMinus_L3D4L4D4_L2_PT_L2L4F2_Minus),
.number_in_projin_layer_10(TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus_number),
.read_add_projin_layer_10(TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus_read_add),
.projin_layer_10(TPROJ_ToMinus_L5D3L6D3_L2_PT_L2L4F2_Minus),
.number_in_projin_layer_11(TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus_number),
.read_add_projin_layer_11(TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus_read_add),
.projin_layer_11(TPROJ_ToMinus_L5D3L6D4_L2_PT_L2L4F2_Minus),
.number_in_projin_layer_12(TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus_number),
.read_add_projin_layer_12(TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus_read_add),
.projin_layer_12(TPROJ_ToMinus_L5D4L6D4_L2_PT_L2L4F2_Minus),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L2L4F2_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L2L4F2_Minus_From_DataStream),
.projout_layer_1(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L3L4),
.valid_layer_1(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L3L4_wr_en),
.projout_layer_2(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L3L4),
.valid_layer_2(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L3L4_wr_en),
.projout_layer_3(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L1L2),
.valid_layer_3(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L1L2_wr_en),
.projout_layer_4(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L1L2),
.valid_layer_4(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L1L2_wr_en),
.projout_layer_5(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L5L6),
.valid_layer_5(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D3_L5L6_wr_en),
.projout_layer_6(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L5L6),
.valid_layer_6(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D3_L5L6_wr_en),
.projout_layer_7(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L5L6),
.valid_layer_7(PT_L2L4F2_Minus_TPROJ_FromMinus_L2D4_L5L6_wr_en),
.projout_layer_8(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L5L6),
.valid_layer_8(PT_L2L4F2_Minus_TPROJ_FromMinus_L4D4_L5L6_wr_en),
.valid_proj_data_stream(PT_L2L4F2_Minus_To_DataStream_en),
.proj_data_stream(PT_L2L4F2_Minus_To_DataStream),
.start(TPROJ_ToMinus_L5D4L6D4_L4_start),
.done(PT_L2L4F2_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("F1L5") PT_F1L5_Minus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus_number),
.read_add_projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus_read_add),
.projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L5_PT_F1L5_Minus),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus_number),
.read_add_projin_layer_4(TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus_read_add),
.projin_layer_4(TPROJ_ToMinus_L3D3L4D3_L5_PT_F1L5_Minus),
.number_in_projin_layer_5(TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus_number),
.read_add_projin_layer_5(TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus_read_add),
.projin_layer_5(TPROJ_ToMinus_L3D3L4D4_L5_PT_F1L5_Minus),
.number_in_projin_layer_6(TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus_number),
.read_add_projin_layer_6(TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus_read_add),
.projin_layer_6(TPROJ_ToMinus_L3D4L4D4_L5_PT_F1L5_Minus),
.number_in_projin_layer_7(6'b0),
.number_in_projin_layer_8(6'b0),
.number_in_projin_layer_9(6'b0),
.number_in_projin_layer_10(6'b0),
.number_in_projin_layer_11(6'b0),
.number_in_projin_layer_12(6'b0),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_F1L5_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_F1L5_Minus_From_DataStream),
.projout_layer_1(PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L3L4),
.valid_layer_1(PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L3L4_wr_en),
.projout_layer_2(PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L3L4),
.valid_layer_2(PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L3L4_wr_en),
.projout_layer_3(PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L1L2),
.valid_layer_3(PT_F1L5_Minus_TPROJ_FromMinus_L5D3_L1L2_wr_en),
.projout_layer_4(PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L1L2),
.valid_layer_4(PT_F1L5_Minus_TPROJ_FromMinus_L5D4_L1L2_wr_en),
.valid_proj_data_stream(PT_F1L5_Minus_To_DataStream_en),
.proj_data_stream(PT_F1L5_Minus_To_DataStream),
.start(TPROJ_ToMinus_L3D4L4D4_L5_start),
.done(PT_F1L5_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionTransceiver #("L1L6F4") PT_L1L6F4_Minus(
.number_in_projin_disk_1(6'b0),
.number_in_projin_disk_2(6'b0),
.number_in_projin_disk_3(6'b0),
.number_in_projin_disk_4(6'b0),
.number_in_projin_disk_5(6'b0),
.number_in_projin_disk_6(6'b0),
.number_in_projin_disk_7(6'b0),
.number_in_projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus_number),
.read_add_projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus_read_add),
.projin_layer_1(TPROJ_ToMinus_L1D3L2D3_L6_PT_L1L6F4_Minus),
.number_in_projin_layer_2(6'b0),
.number_in_projin_layer_3(6'b0),
.number_in_projin_layer_4(TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus_number),
.read_add_projin_layer_4(TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus_read_add),
.projin_layer_4(TPROJ_ToMinus_L3D3L4D3_L6_PT_L1L6F4_Minus),
.number_in_projin_layer_5(TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus_number),
.read_add_projin_layer_5(TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus_read_add),
.projin_layer_5(TPROJ_ToMinus_L3D3L4D4_L6_PT_L1L6F4_Minus),
.number_in_projin_layer_6(TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus_number),
.read_add_projin_layer_6(TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus_read_add),
.projin_layer_6(TPROJ_ToMinus_L3D4L4D4_L6_PT_L1L6F4_Minus),
.number_in_projin_layer_7(TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus_number),
.read_add_projin_layer_7(TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus_read_add),
.projin_layer_7(TPROJ_ToMinus_L3D3L4D3_L1_PT_L1L6F4_Minus),
.number_in_projin_layer_8(TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus_number),
.read_add_projin_layer_8(TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus_read_add),
.projin_layer_8(TPROJ_ToMinus_L3D3L4D4_L1_PT_L1L6F4_Minus),
.number_in_projin_layer_9(TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus_number),
.read_add_projin_layer_9(TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus_read_add),
.projin_layer_9(TPROJ_ToMinus_L3D4L4D4_L1_PT_L1L6F4_Minus),
.number_in_projin_layer_10(TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus_number),
.read_add_projin_layer_10(TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus_read_add),
.projin_layer_10(TPROJ_ToMinus_L5D3L6D3_L1_PT_L1L6F4_Minus),
.number_in_projin_layer_11(TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus_number),
.read_add_projin_layer_11(TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus_read_add),
.projin_layer_11(TPROJ_ToMinus_L5D3L6D4_L1_PT_L1L6F4_Minus),
.number_in_projin_layer_12(TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus_number),
.read_add_projin_layer_12(TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus_read_add),
.projin_layer_12(TPROJ_ToMinus_L5D4L6D4_L1_PT_L1L6F4_Minus),
.number_in_projin_layer_13(6'b0),
.valid_incomming_proj_data_stream(PT_L1L6F4_Minus_From_DataStream_en),
.incomming_proj_data_stream(PT_L1L6F4_Minus_From_DataStream),
.projout_layer_1(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L3L4),
.valid_layer_1(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L3L4_wr_en),
.projout_layer_2(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L3L4),
.valid_layer_2(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L3L4_wr_en),
.projout_layer_3(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L3L4),
.valid_layer_3(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L3L4_wr_en),
.projout_layer_4(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L3L4),
.valid_layer_4(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L3L4_wr_en),
.projout_layer_5(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L1L2),
.valid_layer_5(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D3_L1L2_wr_en),
.projout_layer_6(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L1L2),
.valid_layer_6(PT_L1L6F4_Minus_TPROJ_FromMinus_L6D4_L1L2_wr_en),
.projout_layer_7(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L5L6),
.valid_layer_7(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D3_L5L6_wr_en),
.projout_layer_8(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L5L6),
.valid_layer_8(PT_L1L6F4_Minus_TPROJ_FromMinus_L1D4_L5L6_wr_en),
.valid_proj_data_stream(PT_L1L6F4_Minus_To_DataStream_en),
.proj_data_stream(PT_L1L6F4_Minus_To_DataStream),
.start(TPROJ_ToMinus_L5D4L6D4_L1_start),
.done(PT_L1L6F4_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b1) PR_L1D3_L3L4(
.number_in_proj1in(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_number),
.read_add_proj1in(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L1D3_L3L4_PR_L1D3_L3L4),
.number_in_proj2in(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_number),
.read_add_proj2in(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L1D3_L3L4_PR_L1D3_L3L4),
.number_in_proj3in(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_number),
.read_add_proj3in(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L1D3_PR_L1D3_L3L4),
.number_in_proj4in(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_number),
.read_add_proj4in(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L1D3_PR_L1D3_L3L4),
.number_in_proj5in(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_number),
.read_add_proj5in(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L1D3_PR_L1D3_L3L4),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X1),
.vmprojoutPHI1X2(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X2),
.vmprojoutPHI2X1(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X1),
.vmprojoutPHI2X2(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X2),
.vmprojoutPHI3X1(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X1),
.vmprojoutPHI3X2(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X2),
.allprojout(PR_L1D3_L3L4_AP_L3L4_L1D3),
.valid_data(PR_L1D3_L3L4_AP_L3L4_L1D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L1D3_L3L4_VMPROJ_L3L4_L1D3PHI3X2_wr_en),
.start(TPROJ_FromPlus_L1D3_L3L4_start),
.done(PR_L1D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b1) PR_L2D3_L3L4(
.number_in_proj1in(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_number),
.read_add_proj1in(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L2D3_L3L4_PR_L2D3_L3L4),
.number_in_proj2in(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_number),
.read_add_proj2in(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L2D3_L3L4_PR_L2D3_L3L4),
.number_in_proj3in(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_number),
.read_add_proj3in(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L2D3_PR_L2D3_L3L4),
.number_in_proj4in(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_number),
.read_add_proj4in(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L2D3_PR_L2D3_L3L4),
.number_in_proj5in(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_number),
.read_add_proj5in(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L2D3_PR_L2D3_L3L4),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X1),
.vmprojoutPHI1X2(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X2),
.vmprojoutPHI2X1(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X1),
.vmprojoutPHI2X2(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X2),
.vmprojoutPHI3X1(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X1),
.vmprojoutPHI3X2(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X2),
.vmprojoutPHI4X1(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X1),
.vmprojoutPHI4X2(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X2),
.allprojout(PR_L2D3_L3L4_AP_L3L4_L2D3),
.valid_data(PR_L2D3_L3L4_AP_L3L4_L2D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L2D3_L3L4_VMPROJ_L3L4_L2D3PHI4X2_wr_en),
.start(TPROJ_FromPlus_L2D3_L3L4_start),
.done(PR_L2D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b0) PR_L5D3_L3L4(
.number_in_proj1in(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_number),
.read_add_proj1in(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L5D3_L3L4_PR_L5D3_L3L4),
.number_in_proj2in(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_number),
.read_add_proj2in(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L5D3_L3L4_PR_L5D3_L3L4),
.number_in_proj3in(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_number),
.read_add_proj3in(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L5D3_PR_L5D3_L3L4),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X1),
.vmprojoutPHI1X2(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X2),
.vmprojoutPHI2X1(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X1),
.vmprojoutPHI2X2(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X2),
.vmprojoutPHI3X1(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X1),
.vmprojoutPHI3X2(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X2),
.allprojout(PR_L5D3_L3L4_AP_L3L4_L5D3),
.valid_data(PR_L5D3_L3L4_AP_L3L4_L5D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L5D3_L3L4_VMPROJ_L3L4_L5D3PHI3X2_wr_en),
.start(TPROJ_FromPlus_L5D3_L3L4_start),
.done(PR_L5D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0) PR_L6D3_L3L4(
.number_in_proj1in(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_number),
.read_add_proj1in(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L6D3_L3L4_PR_L6D3_L3L4),
.number_in_proj2in(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_number),
.read_add_proj2in(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L6D3_L3L4_PR_L6D3_L3L4),
.number_in_proj3in(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_number),
.read_add_proj3in(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L6D3_PR_L6D3_L3L4),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X1),
.vmprojoutPHI1X2(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X2),
.vmprojoutPHI2X1(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X1),
.vmprojoutPHI2X2(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X2),
.vmprojoutPHI3X1(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X1),
.vmprojoutPHI3X2(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X2),
.vmprojoutPHI4X1(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X1),
.vmprojoutPHI4X2(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X2),
.allprojout(PR_L6D3_L3L4_AP_L3L4_L6D3),
.valid_data(PR_L6D3_L3L4_AP_L3L4_L6D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L6D3_L3L4_VMPROJ_L3L4_L6D3PHI4X2_wr_en),
.start(TPROJ_FromPlus_L6D3_L3L4_start),
.done(PR_L6D3_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b1) PR_L1D4_L3L4(
.number_in_proj1in(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_number),
.read_add_proj1in(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L1D4_L3L4_PR_L1D4_L3L4),
.number_in_proj2in(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_number),
.read_add_proj2in(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L1D4_L3L4_PR_L1D4_L3L4),
.number_in_proj3in(6'b0),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X1),
.vmprojoutPHI1X2(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X2),
.vmprojoutPHI2X1(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X1),
.vmprojoutPHI2X2(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X2),
.vmprojoutPHI3X1(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X1),
.vmprojoutPHI3X2(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X2),
.allprojout(PR_L1D4_L3L4_AP_L3L4_L1D4),
.valid_data(PR_L1D4_L3L4_AP_L3L4_L1D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L1D4_L3L4_VMPROJ_L3L4_L1D4PHI3X2_wr_en),
.start(TPROJ_FromPlus_L1D4_L3L4_start),
.done(PR_L1D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b1) PR_L2D4_L3L4(
.number_in_proj1in(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_number),
.read_add_proj1in(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L2D4_L3L4_PR_L2D4_L3L4),
.number_in_proj2in(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_number),
.read_add_proj2in(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L2D4_L3L4_PR_L2D4_L3L4),
.number_in_proj3in(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_number),
.read_add_proj3in(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4_read_add),
.proj3in(TPROJ_L3D4L4D4_L2D4_PR_L2D4_L3L4),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X1),
.vmprojoutPHI1X2(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X2),
.vmprojoutPHI2X1(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X1),
.vmprojoutPHI2X2(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X2),
.vmprojoutPHI3X1(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X1),
.vmprojoutPHI3X2(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X2),
.vmprojoutPHI4X1(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X1),
.vmprojoutPHI4X2(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X2),
.allprojout(PR_L2D4_L3L4_AP_L3L4_L2D4),
.valid_data(PR_L2D4_L3L4_AP_L3L4_L2D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L2D4_L3L4_VMPROJ_L3L4_L2D4PHI4X2_wr_en),
.start(TPROJ_FromPlus_L2D4_L3L4_start),
.done(PR_L2D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b0) PR_L5D4_L3L4(
.number_in_proj1in(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_number),
.read_add_proj1in(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L5D4_L3L4_PR_L5D4_L3L4),
.number_in_proj2in(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_number),
.read_add_proj2in(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L5D4_L3L4_PR_L5D4_L3L4),
.number_in_proj3in(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_number),
.read_add_proj3in(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L5D4_PR_L5D4_L3L4),
.number_in_proj4in(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_number),
.read_add_proj4in(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L5D4_PR_L5D4_L3L4),
.number_in_proj5in(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_number),
.read_add_proj5in(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L5D4_PR_L5D4_L3L4),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X1),
.vmprojoutPHI1X2(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X2),
.vmprojoutPHI2X1(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X1),
.vmprojoutPHI2X2(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X2),
.vmprojoutPHI3X1(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X1),
.vmprojoutPHI3X2(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X2),
.allprojout(PR_L5D4_L3L4_AP_L3L4_L5D4),
.valid_data(PR_L5D4_L3L4_AP_L3L4_L5D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L5D4_L3L4_VMPROJ_L3L4_L5D4PHI3X2_wr_en),
.start(TPROJ_FromPlus_L5D4_L3L4_start),
.done(PR_L5D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0) PR_L6D4_L3L4(
.number_in_proj1in(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_number),
.read_add_proj1in(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4_read_add),
.proj1in(TPROJ_FromPlus_L6D4_L3L4_PR_L6D4_L3L4),
.number_in_proj2in(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_number),
.read_add_proj2in(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4_read_add),
.proj2in(TPROJ_FromMinus_L6D4_L3L4_PR_L6D4_L3L4),
.number_in_proj3in(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_number),
.read_add_proj3in(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4_read_add),
.proj3in(TPROJ_L3D3L4D3_L6D4_PR_L6D4_L3L4),
.number_in_proj4in(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_number),
.read_add_proj4in(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4_read_add),
.proj4in(TPROJ_L3D3L4D4_L6D4_PR_L6D4_L3L4),
.number_in_proj5in(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_number),
.read_add_proj5in(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4_read_add),
.proj5in(TPROJ_L3D4L4D4_L6D4_PR_L6D4_L3L4),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X1),
.vmprojoutPHI1X2(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X2),
.vmprojoutPHI2X1(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X1),
.vmprojoutPHI2X2(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X2),
.vmprojoutPHI3X1(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X1),
.vmprojoutPHI3X2(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X2),
.vmprojoutPHI4X1(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X1),
.vmprojoutPHI4X2(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X2),
.allprojout(PR_L6D4_L3L4_AP_L3L4_L6D4),
.valid_data(PR_L6D4_L3L4_AP_L3L4_L6D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L6D4_L3L4_VMPROJ_L3L4_L6D4PHI4X2_wr_en),
.start(TPROJ_FromPlus_L6D4_L3L4_start),
.done(PR_L6D4_L3L4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b1) PR_L3D3_L1L2(
.number_in_proj1in(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_number),
.read_add_proj1in(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L3D3_L1L2_PR_L3D3_L1L2),
.number_in_proj2in(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_number),
.read_add_proj2in(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L3D3_L1L2_PR_L3D3_L1L2),
.number_in_proj3in(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_number),
.read_add_proj3in(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L3D3_PR_L3D3_L1L2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X1),
.vmprojoutPHI1X2(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X2),
.vmprojoutPHI2X1(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X1),
.vmprojoutPHI2X2(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X2),
.vmprojoutPHI3X1(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X1),
.vmprojoutPHI3X2(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X2),
.allprojout(PR_L3D3_L1L2_AP_L1L2_L3D3),
.valid_data(PR_L3D3_L1L2_AP_L1L2_L3D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L3D3_L1L2_VMPROJ_L1L2_L3D3PHI3X2_wr_en),
.start(TPROJ_FromPlus_L3D3_L1L2_start),
.done(PR_L3D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0) PR_L4D3_L1L2(
.number_in_proj1in(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_number),
.read_add_proj1in(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L4D3_L1L2_PR_L4D3_L1L2),
.number_in_proj2in(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_number),
.read_add_proj2in(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L4D3_L1L2_PR_L4D3_L1L2),
.number_in_proj3in(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_number),
.read_add_proj3in(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L4D3_PR_L4D3_L1L2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X1),
.vmprojoutPHI1X2(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X2),
.vmprojoutPHI2X1(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X1),
.vmprojoutPHI2X2(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X2),
.vmprojoutPHI3X1(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X1),
.vmprojoutPHI3X2(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X2),
.vmprojoutPHI4X1(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X1),
.vmprojoutPHI4X2(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X2),
.allprojout(PR_L4D3_L1L2_AP_L1L2_L4D3),
.valid_data(PR_L4D3_L1L2_AP_L1L2_L4D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L4D3_L1L2_VMPROJ_L1L2_L4D3PHI4X2_wr_en),
.start(TPROJ_FromPlus_L4D3_L1L2_start),
.done(PR_L4D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b0) PR_L5D3_L1L2(
.number_in_proj1in(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_number),
.read_add_proj1in(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L5D3_L1L2_PR_L5D3_L1L2),
.number_in_proj2in(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_number),
.read_add_proj2in(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L5D3_L1L2_PR_L5D3_L1L2),
.number_in_proj3in(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_number),
.read_add_proj3in(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L5D3_PR_L5D3_L1L2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X1),
.vmprojoutPHI1X2(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X2),
.vmprojoutPHI2X1(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X1),
.vmprojoutPHI2X2(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X2),
.vmprojoutPHI3X1(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X1),
.vmprojoutPHI3X2(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X2),
.allprojout(PR_L5D3_L1L2_AP_L1L2_L5D3),
.valid_data(PR_L5D3_L1L2_AP_L1L2_L5D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L5D3_L1L2_VMPROJ_L1L2_L5D3PHI3X2_wr_en),
.start(TPROJ_FromPlus_L5D3_L1L2_start),
.done(PR_L5D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0) PR_L6D3_L1L2(
.number_in_proj1in(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_number),
.read_add_proj1in(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L6D3_L1L2_PR_L6D3_L1L2),
.number_in_proj2in(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_number),
.read_add_proj2in(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L6D3_L1L2_PR_L6D3_L1L2),
.number_in_proj3in(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_number),
.read_add_proj3in(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L6D3_PR_L6D3_L1L2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X1),
.vmprojoutPHI1X2(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X2),
.vmprojoutPHI2X1(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X1),
.vmprojoutPHI2X2(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X2),
.vmprojoutPHI3X1(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X1),
.vmprojoutPHI3X2(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X2),
.vmprojoutPHI4X1(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X1),
.vmprojoutPHI4X2(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X2),
.allprojout(PR_L6D3_L1L2_AP_L1L2_L6D3),
.valid_data(PR_L6D3_L1L2_AP_L1L2_L6D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L6D3_L1L2_VMPROJ_L1L2_L6D3PHI4X2_wr_en),
.start(TPROJ_FromPlus_L6D3_L1L2_start),
.done(PR_L6D3_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b1) PR_L3D4_L1L2(
.number_in_proj1in(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_number),
.read_add_proj1in(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L3D4_L1L2_PR_L3D4_L1L2),
.number_in_proj2in(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_number),
.read_add_proj2in(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L3D4_L1L2_PR_L3D4_L1L2),
.number_in_proj3in(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_number),
.read_add_proj3in(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L3D4_PR_L3D4_L1L2),
.number_in_proj4in(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_number),
.read_add_proj4in(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L3D4_PR_L3D4_L1L2),
.number_in_proj5in(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_number),
.read_add_proj5in(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2_read_add),
.proj5in(TPROJ_L1D4L2D4_L3D4_PR_L3D4_L1L2),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X1),
.vmprojoutPHI1X2(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X2),
.vmprojoutPHI2X1(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X1),
.vmprojoutPHI2X2(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X2),
.vmprojoutPHI3X1(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X1),
.vmprojoutPHI3X2(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X2),
.allprojout(PR_L3D4_L1L2_AP_L1L2_L3D4),
.valid_data(PR_L3D4_L1L2_AP_L1L2_L3D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L3D4_L1L2_VMPROJ_L1L2_L3D4PHI3X2_wr_en),
.start(TPROJ_FromPlus_L3D4_L1L2_start),
.done(PR_L3D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0) PR_L4D4_L1L2(
.number_in_proj1in(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_number),
.read_add_proj1in(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L4D4_L1L2_PR_L4D4_L1L2),
.number_in_proj2in(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_number),
.read_add_proj2in(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L4D4_L1L2_PR_L4D4_L1L2),
.number_in_proj3in(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_number),
.read_add_proj3in(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L4D4_PR_L4D4_L1L2),
.number_in_proj4in(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_number),
.read_add_proj4in(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2_read_add),
.proj4in(TPROJ_L1D3L2D4_L4D4_PR_L4D4_L1L2),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X1),
.vmprojoutPHI1X2(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X2),
.vmprojoutPHI2X1(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X1),
.vmprojoutPHI2X2(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X2),
.vmprojoutPHI3X1(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X1),
.vmprojoutPHI3X2(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X2),
.vmprojoutPHI4X1(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X1),
.vmprojoutPHI4X2(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X2),
.allprojout(PR_L4D4_L1L2_AP_L1L2_L4D4),
.valid_data(PR_L4D4_L1L2_AP_L1L2_L4D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L4D4_L1L2_VMPROJ_L1L2_L4D4PHI4X2_wr_en),
.start(TPROJ_FromPlus_L4D4_L1L2_start),
.done(PR_L4D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b0) PR_L5D4_L1L2(
.number_in_proj1in(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_number),
.read_add_proj1in(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L5D4_L1L2_PR_L5D4_L1L2),
.number_in_proj2in(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_number),
.read_add_proj2in(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L5D4_L1L2_PR_L5D4_L1L2),
.number_in_proj3in(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_number),
.read_add_proj3in(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L5D4_PR_L5D4_L1L2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X1),
.vmprojoutPHI1X2(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X2),
.vmprojoutPHI2X1(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X1),
.vmprojoutPHI2X2(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X2),
.vmprojoutPHI3X1(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X1),
.vmprojoutPHI3X2(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X2),
.allprojout(PR_L5D4_L1L2_AP_L1L2_L5D4),
.valid_data(PR_L5D4_L1L2_AP_L1L2_L5D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L5D4_L1L2_VMPROJ_L1L2_L5D4PHI3X2_wr_en),
.start(TPROJ_FromPlus_L5D4_L1L2_start),
.done(PR_L5D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0) PR_L6D4_L1L2(
.number_in_proj1in(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_number),
.read_add_proj1in(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2_read_add),
.proj1in(TPROJ_FromPlus_L6D4_L1L2_PR_L6D4_L1L2),
.number_in_proj2in(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_number),
.read_add_proj2in(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2_read_add),
.proj2in(TPROJ_FromMinus_L6D4_L1L2_PR_L6D4_L1L2),
.number_in_proj3in(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_number),
.read_add_proj3in(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2_read_add),
.proj3in(TPROJ_L1D3L2D3_L6D4_PR_L6D4_L1L2),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X1),
.vmprojoutPHI1X2(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X2),
.vmprojoutPHI2X1(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X1),
.vmprojoutPHI2X2(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X2),
.vmprojoutPHI3X1(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X1),
.vmprojoutPHI3X2(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X2),
.vmprojoutPHI4X1(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X1),
.vmprojoutPHI4X2(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X2),
.allprojout(PR_L6D4_L1L2_AP_L1L2_L6D4),
.valid_data(PR_L6D4_L1L2_AP_L1L2_L6D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L6D4_L1L2_VMPROJ_L1L2_L6D4PHI4X2_wr_en),
.start(TPROJ_FromPlus_L6D4_L1L2_start),
.done(PR_L6D4_L1L2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b1) PR_L1D3_L5L6(
.number_in_proj1in(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_number),
.read_add_proj1in(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L1D3_L5L6_PR_L1D3_L5L6),
.number_in_proj2in(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_number),
.read_add_proj2in(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L1D3_L5L6_PR_L1D3_L5L6),
.number_in_proj3in(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_number),
.read_add_proj3in(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L1D3_PR_L1D3_L5L6),
.number_in_proj4in(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_number),
.read_add_proj4in(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L1D3_PR_L1D3_L5L6),
.number_in_proj5in(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_number),
.read_add_proj5in(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L1D3_PR_L1D3_L5L6),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X1),
.vmprojoutPHI1X2(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X2),
.vmprojoutPHI2X1(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X1),
.vmprojoutPHI2X2(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X2),
.vmprojoutPHI3X1(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X1),
.vmprojoutPHI3X2(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X2),
.allprojout(PR_L1D3_L5L6_AP_L5L6_L1D3),
.valid_data(PR_L1D3_L5L6_AP_L5L6_L1D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L1D3_L5L6_VMPROJ_L5L6_L1D3PHI3X2_wr_en),
.start(TPROJ_FromPlus_L1D3_L5L6_start),
.done(PR_L1D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b1) PR_L2D3_L5L6(
.number_in_proj1in(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_number),
.read_add_proj1in(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L2D3_L5L6_PR_L2D3_L5L6),
.number_in_proj2in(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_number),
.read_add_proj2in(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L2D3_L5L6_PR_L2D3_L5L6),
.number_in_proj3in(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_number),
.read_add_proj3in(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L2D3_PR_L2D3_L5L6),
.number_in_proj4in(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_number),
.read_add_proj4in(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L2D3_PR_L2D3_L5L6),
.number_in_proj5in(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_number),
.read_add_proj5in(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L2D3_PR_L2D3_L5L6),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X1),
.vmprojoutPHI1X2(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X2),
.vmprojoutPHI2X1(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X1),
.vmprojoutPHI2X2(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X2),
.vmprojoutPHI3X1(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X1),
.vmprojoutPHI3X2(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X2),
.vmprojoutPHI4X1(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X1),
.vmprojoutPHI4X2(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X2),
.allprojout(PR_L2D3_L5L6_AP_L5L6_L2D3),
.valid_data(PR_L2D3_L5L6_AP_L5L6_L2D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L2D3_L5L6_VMPROJ_L5L6_L2D3PHI4X2_wr_en),
.start(TPROJ_FromPlus_L2D3_L5L6_start),
.done(PR_L2D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b1) PR_L3D3_L5L6(
.number_in_proj1in(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_number),
.read_add_proj1in(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L3D3_L5L6_PR_L3D3_L5L6),
.number_in_proj2in(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_number),
.read_add_proj2in(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L3D3_L5L6_PR_L3D3_L5L6),
.number_in_proj3in(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_number),
.read_add_proj3in(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L3D3_PR_L3D3_L5L6),
.number_in_proj4in(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_number),
.read_add_proj4in(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L3D3_PR_L3D3_L5L6),
.number_in_proj5in(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_number),
.read_add_proj5in(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L3D3_PR_L3D3_L5L6),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X1),
.vmprojoutPHI1X2(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X2),
.vmprojoutPHI2X1(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X1),
.vmprojoutPHI2X2(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X2),
.vmprojoutPHI3X1(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X1),
.vmprojoutPHI3X2(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X2),
.allprojout(PR_L3D3_L5L6_AP_L5L6_L3D3),
.valid_data(PR_L3D3_L5L6_AP_L5L6_L3D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L3D3_L5L6_VMPROJ_L5L6_L3D3PHI3X2_wr_en),
.start(TPROJ_FromPlus_L3D3_L5L6_start),
.done(PR_L3D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0) PR_L4D3_L5L6(
.number_in_proj1in(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_number),
.read_add_proj1in(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L4D3_L5L6_PR_L4D3_L5L6),
.number_in_proj2in(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_number),
.read_add_proj2in(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L4D3_L5L6_PR_L4D3_L5L6),
.number_in_proj3in(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_number),
.read_add_proj3in(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6_read_add),
.proj3in(TPROJ_L5D3L6D3_L4D3_PR_L4D3_L5L6),
.number_in_proj4in(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_number),
.read_add_proj4in(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6_read_add),
.proj4in(TPROJ_L5D3L6D4_L4D3_PR_L4D3_L5L6),
.number_in_proj5in(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_number),
.read_add_proj5in(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6_read_add),
.proj5in(TPROJ_L5D4L6D4_L4D3_PR_L4D3_L5L6),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X1),
.vmprojoutPHI1X2(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X2),
.vmprojoutPHI2X1(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X1),
.vmprojoutPHI2X2(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X2),
.vmprojoutPHI3X1(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X1),
.vmprojoutPHI3X2(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X2),
.vmprojoutPHI4X1(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X1),
.vmprojoutPHI4X2(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X2),
.allprojout(PR_L4D3_L5L6_AP_L5L6_L4D3),
.valid_data(PR_L4D3_L5L6_AP_L5L6_L4D3_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L4D3_L5L6_VMPROJ_L5L6_L4D3PHI4X2_wr_en),
.start(TPROJ_FromPlus_L4D3_L5L6_start),
.done(PR_L4D3_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b1) PR_L1D4_L5L6(
.number_in_proj1in(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_number),
.read_add_proj1in(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L1D4_L5L6_PR_L1D4_L5L6),
.number_in_proj2in(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_number),
.read_add_proj2in(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L1D4_L5L6_PR_L1D4_L5L6),
.number_in_proj3in(6'b0),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X1),
.vmprojoutPHI1X2(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X2),
.vmprojoutPHI2X1(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X1),
.vmprojoutPHI2X2(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X2),
.vmprojoutPHI3X1(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X1),
.vmprojoutPHI3X2(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X2),
.allprojout(PR_L1D4_L5L6_AP_L5L6_L1D4),
.valid_data(PR_L1D4_L5L6_AP_L5L6_L1D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L1D4_L5L6_VMPROJ_L5L6_L1D4PHI3X2_wr_en),
.start(TPROJ_FromPlus_L1D4_L5L6_start),
.done(PR_L1D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b1) PR_L2D4_L5L6(
.number_in_proj1in(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_number),
.read_add_proj1in(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L2D4_L5L6_PR_L2D4_L5L6),
.number_in_proj2in(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_number),
.read_add_proj2in(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L2D4_L5L6_PR_L2D4_L5L6),
.number_in_proj3in(6'b0),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X1),
.vmprojoutPHI1X2(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X2),
.vmprojoutPHI2X1(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X1),
.vmprojoutPHI2X2(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X2),
.vmprojoutPHI3X1(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X1),
.vmprojoutPHI3X2(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X2),
.vmprojoutPHI4X1(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X1),
.vmprojoutPHI4X2(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X2),
.allprojout(PR_L2D4_L5L6_AP_L5L6_L2D4),
.valid_data(PR_L2D4_L5L6_AP_L5L6_L2D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L2D4_L5L6_VMPROJ_L5L6_L2D4PHI4X2_wr_en),
.start(TPROJ_FromPlus_L2D4_L5L6_start),
.done(PR_L2D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b1,1'b1) PR_L3D4_L5L6(
.number_in_proj1in(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_number),
.read_add_proj1in(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L3D4_L5L6_PR_L3D4_L5L6),
.number_in_proj2in(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_number),
.read_add_proj2in(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L3D4_L5L6_PR_L3D4_L5L6),
.number_in_proj3in(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_number),
.read_add_proj3in(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6_read_add),
.proj3in(TPROJ_L5D4L6D4_L3D4_PR_L3D4_L5L6),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X1),
.vmprojoutPHI1X2(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X2),
.vmprojoutPHI2X1(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X1),
.vmprojoutPHI2X2(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X2),
.vmprojoutPHI3X1(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X1),
.vmprojoutPHI3X2(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X2),
.allprojout(PR_L3D4_L5L6_AP_L5L6_L3D4),
.valid_data(PR_L3D4_L5L6_AP_L5L6_L3D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L3D4_L5L6_VMPROJ_L5L6_L3D4PHI3X2_wr_en),
.start(TPROJ_FromPlus_L3D4_L5L6_start),
.done(PR_L3D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

ProjectionRouter #(1'b0,1'b0) PR_L4D4_L5L6(
.number_in_proj1in(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_number),
.read_add_proj1in(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6_read_add),
.proj1in(TPROJ_FromPlus_L4D4_L5L6_PR_L4D4_L5L6),
.number_in_proj2in(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_number),
.read_add_proj2in(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6_read_add),
.proj2in(TPROJ_FromMinus_L4D4_L5L6_PR_L4D4_L5L6),
.number_in_proj3in(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_number),
.read_add_proj3in(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6_read_add),
.proj3in(TPROJ_L5D4L6D4_L4D4_PR_L4D4_L5L6),
.number_in_proj4in(6'b0),
.number_in_proj5in(6'b0),
.number_in_proj6in(6'b0),
.number_in_proj7in(6'b0),
.vmprojoutPHI1X1(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X1),
.vmprojoutPHI1X2(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X2),
.vmprojoutPHI2X1(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X1),
.vmprojoutPHI2X2(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X2),
.vmprojoutPHI3X1(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X1),
.vmprojoutPHI3X2(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X2),
.vmprojoutPHI4X1(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X1),
.vmprojoutPHI4X2(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X2),
.allprojout(PR_L4D4_L5L6_AP_L5L6_L4D4),
.valid_data(PR_L4D4_L5L6_AP_L5L6_L4D4_wr_en),
.vmprojoutPHI1X1_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X1_wr_en),
.vmprojoutPHI1X2_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI1X2_wr_en),
.vmprojoutPHI2X1_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X1_wr_en),
.vmprojoutPHI2X2_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI2X2_wr_en),
.vmprojoutPHI3X1_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X1_wr_en),
.vmprojoutPHI3X2_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI3X2_wr_en),
.vmprojoutPHI4X1_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X1_wr_en),
.vmprojoutPHI4X2_wr_en(PR_L4D4_L5L6_VMPROJ_L5L6_L4D4PHI4X2_wr_en),
.start(TPROJ_FromPlus_L4D4_L5L6_start),
.done(PR_L4D4_L5L6_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D3PHI1X1(
.number_in_vmstubin(VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1_number),
.read_add_vmstubin(VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1_read_add),
.vmstubin(VMS_L1D3PHI1X1n7_ME_L3L4_L1D3PHI1X1),
.number_in_vmprojin(VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI1X1_ME_L3L4_L1D3PHI1X1),
.matchout(ME_L3L4_L1D3PHI1X1_CM_L3L4_L1D3PHI1X1),
.valid_data(ME_L3L4_L1D3PHI1X1_CM_L3L4_L1D3PHI1X1_wr_en),
.start(VMPROJ_L3L4_L1D3PHI1X1_start),
.done(ME_L3L4_L1D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D3PHI1X2(
.number_in_vmstubin(VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2_number),
.read_add_vmstubin(VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2_read_add),
.vmstubin(VMS_L1D3PHI1X2n7_ME_L3L4_L1D3PHI1X2),
.number_in_vmprojin(VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI1X2_ME_L3L4_L1D3PHI1X2),
.matchout(ME_L3L4_L1D3PHI1X2_CM_L3L4_L1D3PHI1X2),
.valid_data(ME_L3L4_L1D3PHI1X2_CM_L3L4_L1D3PHI1X2_wr_en),
.start(VMPROJ_L3L4_L1D3PHI1X2_start),
.done(ME_L3L4_L1D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D3PHI2X1(
.number_in_vmstubin(VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1_number),
.read_add_vmstubin(VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1_read_add),
.vmstubin(VMS_L1D3PHI2X1n7_ME_L3L4_L1D3PHI2X1),
.number_in_vmprojin(VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI2X1_ME_L3L4_L1D3PHI2X1),
.matchout(ME_L3L4_L1D3PHI2X1_CM_L3L4_L1D3PHI2X1),
.valid_data(ME_L3L4_L1D3PHI2X1_CM_L3L4_L1D3PHI2X1_wr_en),
.start(VMPROJ_L3L4_L1D3PHI2X1_start),
.done(ME_L3L4_L1D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D3PHI2X2(
.number_in_vmstubin(VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2_number),
.read_add_vmstubin(VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2_read_add),
.vmstubin(VMS_L1D3PHI2X2n7_ME_L3L4_L1D3PHI2X2),
.number_in_vmprojin(VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI2X2_ME_L3L4_L1D3PHI2X2),
.matchout(ME_L3L4_L1D3PHI2X2_CM_L3L4_L1D3PHI2X2),
.valid_data(ME_L3L4_L1D3PHI2X2_CM_L3L4_L1D3PHI2X2_wr_en),
.start(VMPROJ_L3L4_L1D3PHI2X2_start),
.done(ME_L3L4_L1D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D3PHI3X1(
.number_in_vmstubin(VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1_number),
.read_add_vmstubin(VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1_read_add),
.vmstubin(VMS_L1D3PHI3X1n7_ME_L3L4_L1D3PHI3X1),
.number_in_vmprojin(VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI3X1_ME_L3L4_L1D3PHI3X1),
.matchout(ME_L3L4_L1D3PHI3X1_CM_L3L4_L1D3PHI3X1),
.valid_data(ME_L3L4_L1D3PHI3X1_CM_L3L4_L1D3PHI3X1_wr_en),
.start(VMPROJ_L3L4_L1D3PHI3X1_start),
.done(ME_L3L4_L1D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D3PHI3X2(
.number_in_vmstubin(VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2_number),
.read_add_vmstubin(VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2_read_add),
.vmstubin(VMS_L1D3PHI3X2n7_ME_L3L4_L1D3PHI3X2),
.number_in_vmprojin(VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2_read_add),
.vmprojin(VMPROJ_L3L4_L1D3PHI3X2_ME_L3L4_L1D3PHI3X2),
.matchout(ME_L3L4_L1D3PHI3X2_CM_L3L4_L1D3PHI3X2),
.valid_data(ME_L3L4_L1D3PHI3X2_CM_L3L4_L1D3PHI3X2_wr_en),
.start(VMPROJ_L3L4_L1D3PHI3X2_start),
.done(ME_L3L4_L1D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D4PHI1X1(
.number_in_vmstubin(VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1_number),
.read_add_vmstubin(VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1_read_add),
.vmstubin(VMS_L1D4PHI1X1n3_ME_L3L4_L1D4PHI1X1),
.number_in_vmprojin(VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI1X1_ME_L3L4_L1D4PHI1X1),
.matchout(ME_L3L4_L1D4PHI1X1_CM_L3L4_L1D4PHI1X1),
.valid_data(ME_L3L4_L1D4PHI1X1_CM_L3L4_L1D4PHI1X1_wr_en),
.start(VMPROJ_L3L4_L1D4PHI1X1_start),
.done(ME_L3L4_L1D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D4PHI1X2(
.number_in_vmprojin(VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI1X2_ME_L3L4_L1D4PHI1X2),
.number_in_vmstubin(VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2_number),
.read_add_vmstubin(VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2_read_add),
.vmstubin(VMS_L1D4PHI1X2n1_ME_L3L4_L1D4PHI1X2),
.matchout(ME_L3L4_L1D4PHI1X2_CM_L3L4_L1D4PHI1X2),
.valid_data(ME_L3L4_L1D4PHI1X2_CM_L3L4_L1D4PHI1X2_wr_en),
.start(VMPROJ_L3L4_L1D4PHI1X2_start),
.done(ME_L3L4_L1D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D4PHI2X1(
.number_in_vmstubin(VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1_number),
.read_add_vmstubin(VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1_read_add),
.vmstubin(VMS_L1D4PHI2X1n3_ME_L3L4_L1D4PHI2X1),
.number_in_vmprojin(VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI2X1_ME_L3L4_L1D4PHI2X1),
.matchout(ME_L3L4_L1D4PHI2X1_CM_L3L4_L1D4PHI2X1),
.valid_data(ME_L3L4_L1D4PHI2X1_CM_L3L4_L1D4PHI2X1_wr_en),
.start(VMPROJ_L3L4_L1D4PHI2X1_start),
.done(ME_L3L4_L1D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D4PHI2X2(
.number_in_vmprojin(VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI2X2_ME_L3L4_L1D4PHI2X2),
.number_in_vmstubin(VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2_number),
.read_add_vmstubin(VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2_read_add),
.vmstubin(VMS_L1D4PHI2X2n1_ME_L3L4_L1D4PHI2X2),
.matchout(ME_L3L4_L1D4PHI2X2_CM_L3L4_L1D4PHI2X2),
.valid_data(ME_L3L4_L1D4PHI2X2_CM_L3L4_L1D4PHI2X2_wr_en),
.start(VMPROJ_L3L4_L1D4PHI2X2_start),
.done(ME_L3L4_L1D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D4PHI3X1(
.number_in_vmstubin(VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1_number),
.read_add_vmstubin(VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1_read_add),
.vmstubin(VMS_L1D4PHI3X1n3_ME_L3L4_L1D4PHI3X1),
.number_in_vmprojin(VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI3X1_ME_L3L4_L1D4PHI3X1),
.matchout(ME_L3L4_L1D4PHI3X1_CM_L3L4_L1D4PHI3X1),
.valid_data(ME_L3L4_L1D4PHI3X1_CM_L3L4_L1D4PHI3X1_wr_en),
.start(VMPROJ_L3L4_L1D4PHI3X1_start),
.done(ME_L3L4_L1D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L1D4PHI3X2(
.number_in_vmprojin(VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2_read_add),
.vmprojin(VMPROJ_L3L4_L1D4PHI3X2_ME_L3L4_L1D4PHI3X2),
.number_in_vmstubin(VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2_number),
.read_add_vmstubin(VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2_read_add),
.vmstubin(VMS_L1D4PHI3X2n1_ME_L3L4_L1D4PHI3X2),
.matchout(ME_L3L4_L1D4PHI3X2_CM_L3L4_L1D4PHI3X2),
.valid_data(ME_L3L4_L1D4PHI3X2_CM_L3L4_L1D4PHI3X2_wr_en),
.start(VMPROJ_L3L4_L1D4PHI3X2_start),
.done(ME_L3L4_L1D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D3PHI1X1(
.number_in_vmstubin(VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1_number),
.read_add_vmstubin(VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1_read_add),
.vmstubin(VMS_L2D3PHI1X1n2_ME_L3L4_L2D3PHI1X1),
.number_in_vmprojin(VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI1X1_ME_L3L4_L2D3PHI1X1),
.matchout(ME_L3L4_L2D3PHI1X1_CM_L3L4_L2D3PHI1X1),
.valid_data(ME_L3L4_L2D3PHI1X1_CM_L3L4_L2D3PHI1X1_wr_en),
.start(VMPROJ_L3L4_L2D3PHI1X1_start),
.done(ME_L3L4_L2D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D3PHI1X2(
.number_in_vmstubin(VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2_number),
.read_add_vmstubin(VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2_read_add),
.vmstubin(VMS_L2D3PHI1X2n3_ME_L3L4_L2D3PHI1X2),
.number_in_vmprojin(VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI1X2_ME_L3L4_L2D3PHI1X2),
.matchout(ME_L3L4_L2D3PHI1X2_CM_L3L4_L2D3PHI1X2),
.valid_data(ME_L3L4_L2D3PHI1X2_CM_L3L4_L2D3PHI1X2_wr_en),
.start(VMPROJ_L3L4_L2D3PHI1X2_start),
.done(ME_L3L4_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D3PHI2X1(
.number_in_vmstubin(VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1_number),
.read_add_vmstubin(VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1_read_add),
.vmstubin(VMS_L2D3PHI2X1n3_ME_L3L4_L2D3PHI2X1),
.number_in_vmprojin(VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI2X1_ME_L3L4_L2D3PHI2X1),
.matchout(ME_L3L4_L2D3PHI2X1_CM_L3L4_L2D3PHI2X1),
.valid_data(ME_L3L4_L2D3PHI2X1_CM_L3L4_L2D3PHI2X1_wr_en),
.start(VMPROJ_L3L4_L2D3PHI2X1_start),
.done(ME_L3L4_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D3PHI2X2(
.number_in_vmstubin(VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2_number),
.read_add_vmstubin(VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2_read_add),
.vmstubin(VMS_L2D3PHI2X2n5_ME_L3L4_L2D3PHI2X2),
.number_in_vmprojin(VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI2X2_ME_L3L4_L2D3PHI2X2),
.matchout(ME_L3L4_L2D3PHI2X2_CM_L3L4_L2D3PHI2X2),
.valid_data(ME_L3L4_L2D3PHI2X2_CM_L3L4_L2D3PHI2X2_wr_en),
.start(VMPROJ_L3L4_L2D3PHI2X2_start),
.done(ME_L3L4_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D3PHI3X1(
.number_in_vmstubin(VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1_number),
.read_add_vmstubin(VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1_read_add),
.vmstubin(VMS_L2D3PHI3X1n3_ME_L3L4_L2D3PHI3X1),
.number_in_vmprojin(VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI3X1_ME_L3L4_L2D3PHI3X1),
.matchout(ME_L3L4_L2D3PHI3X1_CM_L3L4_L2D3PHI3X1),
.valid_data(ME_L3L4_L2D3PHI3X1_CM_L3L4_L2D3PHI3X1_wr_en),
.start(VMPROJ_L3L4_L2D3PHI3X1_start),
.done(ME_L3L4_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D3PHI3X2(
.number_in_vmstubin(VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2_number),
.read_add_vmstubin(VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2_read_add),
.vmstubin(VMS_L2D3PHI3X2n5_ME_L3L4_L2D3PHI3X2),
.number_in_vmprojin(VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI3X2_ME_L3L4_L2D3PHI3X2),
.matchout(ME_L3L4_L2D3PHI3X2_CM_L3L4_L2D3PHI3X2),
.valid_data(ME_L3L4_L2D3PHI3X2_CM_L3L4_L2D3PHI3X2_wr_en),
.start(VMPROJ_L3L4_L2D3PHI3X2_start),
.done(ME_L3L4_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D3PHI4X1(
.number_in_vmstubin(VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1_number),
.read_add_vmstubin(VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1_read_add),
.vmstubin(VMS_L2D3PHI4X1n2_ME_L3L4_L2D3PHI4X1),
.number_in_vmprojin(VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI4X1_ME_L3L4_L2D3PHI4X1),
.matchout(ME_L3L4_L2D3PHI4X1_CM_L3L4_L2D3PHI4X1),
.valid_data(ME_L3L4_L2D3PHI4X1_CM_L3L4_L2D3PHI4X1_wr_en),
.start(VMPROJ_L3L4_L2D3PHI4X1_start),
.done(ME_L3L4_L2D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D3PHI4X2(
.number_in_vmstubin(VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2_number),
.read_add_vmstubin(VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2_read_add),
.vmstubin(VMS_L2D3PHI4X2n3_ME_L3L4_L2D3PHI4X2),
.number_in_vmprojin(VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2_read_add),
.vmprojin(VMPROJ_L3L4_L2D3PHI4X2_ME_L3L4_L2D3PHI4X2),
.matchout(ME_L3L4_L2D3PHI4X2_CM_L3L4_L2D3PHI4X2),
.valid_data(ME_L3L4_L2D3PHI4X2_CM_L3L4_L2D3PHI4X2_wr_en),
.start(VMPROJ_L3L4_L2D3PHI4X2_start),
.done(ME_L3L4_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D4PHI1X1(
.number_in_vmstubin(VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1_number),
.read_add_vmstubin(VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1_read_add),
.vmstubin(VMS_L2D4PHI1X1n3_ME_L3L4_L2D4PHI1X1),
.number_in_vmprojin(VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI1X1_ME_L3L4_L2D4PHI1X1),
.matchout(ME_L3L4_L2D4PHI1X1_CM_L3L4_L2D4PHI1X1),
.valid_data(ME_L3L4_L2D4PHI1X1_CM_L3L4_L2D4PHI1X1_wr_en),
.start(VMPROJ_L3L4_L2D4PHI1X1_start),
.done(ME_L3L4_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D4PHI1X2(
.number_in_vmstubin(VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2_number),
.read_add_vmstubin(VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2_read_add),
.vmstubin(VMS_L2D4PHI1X2n3_ME_L3L4_L2D4PHI1X2),
.number_in_vmprojin(VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI1X2_ME_L3L4_L2D4PHI1X2),
.matchout(ME_L3L4_L2D4PHI1X2_CM_L3L4_L2D4PHI1X2),
.valid_data(ME_L3L4_L2D4PHI1X2_CM_L3L4_L2D4PHI1X2_wr_en),
.start(VMPROJ_L3L4_L2D4PHI1X2_start),
.done(ME_L3L4_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D4PHI2X1(
.number_in_vmstubin(VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1_number),
.read_add_vmstubin(VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1_read_add),
.vmstubin(VMS_L2D4PHI2X1n5_ME_L3L4_L2D4PHI2X1),
.number_in_vmprojin(VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI2X1_ME_L3L4_L2D4PHI2X1),
.matchout(ME_L3L4_L2D4PHI2X1_CM_L3L4_L2D4PHI2X1),
.valid_data(ME_L3L4_L2D4PHI2X1_CM_L3L4_L2D4PHI2X1_wr_en),
.start(VMPROJ_L3L4_L2D4PHI2X1_start),
.done(ME_L3L4_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D4PHI2X2(
.number_in_vmstubin(VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2_number),
.read_add_vmstubin(VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2_read_add),
.vmstubin(VMS_L2D4PHI2X2n5_ME_L3L4_L2D4PHI2X2),
.number_in_vmprojin(VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI2X2_ME_L3L4_L2D4PHI2X2),
.matchout(ME_L3L4_L2D4PHI2X2_CM_L3L4_L2D4PHI2X2),
.valid_data(ME_L3L4_L2D4PHI2X2_CM_L3L4_L2D4PHI2X2_wr_en),
.start(VMPROJ_L3L4_L2D4PHI2X2_start),
.done(ME_L3L4_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D4PHI3X1(
.number_in_vmstubin(VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1_number),
.read_add_vmstubin(VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1_read_add),
.vmstubin(VMS_L2D4PHI3X1n5_ME_L3L4_L2D4PHI3X1),
.number_in_vmprojin(VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI3X1_ME_L3L4_L2D4PHI3X1),
.matchout(ME_L3L4_L2D4PHI3X1_CM_L3L4_L2D4PHI3X1),
.valid_data(ME_L3L4_L2D4PHI3X1_CM_L3L4_L2D4PHI3X1_wr_en),
.start(VMPROJ_L3L4_L2D4PHI3X1_start),
.done(ME_L3L4_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D4PHI3X2(
.number_in_vmstubin(VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2_number),
.read_add_vmstubin(VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2_read_add),
.vmstubin(VMS_L2D4PHI3X2n5_ME_L3L4_L2D4PHI3X2),
.number_in_vmprojin(VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI3X2_ME_L3L4_L2D4PHI3X2),
.matchout(ME_L3L4_L2D4PHI3X2_CM_L3L4_L2D4PHI3X2),
.valid_data(ME_L3L4_L2D4PHI3X2_CM_L3L4_L2D4PHI3X2_wr_en),
.start(VMPROJ_L3L4_L2D4PHI3X2_start),
.done(ME_L3L4_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D4PHI4X1(
.number_in_vmstubin(VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1_number),
.read_add_vmstubin(VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1_read_add),
.vmstubin(VMS_L2D4PHI4X1n3_ME_L3L4_L2D4PHI4X1),
.number_in_vmprojin(VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI4X1_ME_L3L4_L2D4PHI4X1),
.matchout(ME_L3L4_L2D4PHI4X1_CM_L3L4_L2D4PHI4X1),
.valid_data(ME_L3L4_L2D4PHI4X1_CM_L3L4_L2D4PHI4X1_wr_en),
.start(VMPROJ_L3L4_L2D4PHI4X1_start),
.done(ME_L3L4_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L2D4PHI4X2(
.number_in_vmstubin(VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2_number),
.read_add_vmstubin(VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2_read_add),
.vmstubin(VMS_L2D4PHI4X2n3_ME_L3L4_L2D4PHI4X2),
.number_in_vmprojin(VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2_read_add),
.vmprojin(VMPROJ_L3L4_L2D4PHI4X2_ME_L3L4_L2D4PHI4X2),
.matchout(ME_L3L4_L2D4PHI4X2_CM_L3L4_L2D4PHI4X2),
.valid_data(ME_L3L4_L2D4PHI4X2_CM_L3L4_L2D4PHI4X2_wr_en),
.start(VMPROJ_L3L4_L2D4PHI4X2_start),
.done(ME_L3L4_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D3PHI1X1(
.number_in_vmstubin(VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1_number),
.read_add_vmstubin(VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1_read_add),
.vmstubin(VMS_L5D3PHI1X1n5_ME_L3L4_L5D3PHI1X1),
.number_in_vmprojin(VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI1X1_ME_L3L4_L5D3PHI1X1),
.matchout(ME_L3L4_L5D3PHI1X1_CM_L3L4_L5D3PHI1X1),
.valid_data(ME_L3L4_L5D3PHI1X1_CM_L3L4_L5D3PHI1X1_wr_en),
.start(VMPROJ_L3L4_L5D3PHI1X1_start),
.done(ME_L3L4_L5D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D3PHI1X2(
.number_in_vmstubin(VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2_number),
.read_add_vmstubin(VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2_read_add),
.vmstubin(VMS_L5D3PHI1X2n5_ME_L3L4_L5D3PHI1X2),
.number_in_vmprojin(VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI1X2_ME_L3L4_L5D3PHI1X2),
.matchout(ME_L3L4_L5D3PHI1X2_CM_L3L4_L5D3PHI1X2),
.valid_data(ME_L3L4_L5D3PHI1X2_CM_L3L4_L5D3PHI1X2_wr_en),
.start(VMPROJ_L3L4_L5D3PHI1X2_start),
.done(ME_L3L4_L5D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D3PHI2X1(
.number_in_vmstubin(VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1_number),
.read_add_vmstubin(VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1_read_add),
.vmstubin(VMS_L5D3PHI2X1n5_ME_L3L4_L5D3PHI2X1),
.number_in_vmprojin(VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI2X1_ME_L3L4_L5D3PHI2X1),
.matchout(ME_L3L4_L5D3PHI2X1_CM_L3L4_L5D3PHI2X1),
.valid_data(ME_L3L4_L5D3PHI2X1_CM_L3L4_L5D3PHI2X1_wr_en),
.start(VMPROJ_L3L4_L5D3PHI2X1_start),
.done(ME_L3L4_L5D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D3PHI2X2(
.number_in_vmstubin(VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2_number),
.read_add_vmstubin(VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2_read_add),
.vmstubin(VMS_L5D3PHI2X2n5_ME_L3L4_L5D3PHI2X2),
.number_in_vmprojin(VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI2X2_ME_L3L4_L5D3PHI2X2),
.matchout(ME_L3L4_L5D3PHI2X2_CM_L3L4_L5D3PHI2X2),
.valid_data(ME_L3L4_L5D3PHI2X2_CM_L3L4_L5D3PHI2X2_wr_en),
.start(VMPROJ_L3L4_L5D3PHI2X2_start),
.done(ME_L3L4_L5D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D3PHI3X1(
.number_in_vmstubin(VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1_number),
.read_add_vmstubin(VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1_read_add),
.vmstubin(VMS_L5D3PHI3X1n5_ME_L3L4_L5D3PHI3X1),
.number_in_vmprojin(VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI3X1_ME_L3L4_L5D3PHI3X1),
.matchout(ME_L3L4_L5D3PHI3X1_CM_L3L4_L5D3PHI3X1),
.valid_data(ME_L3L4_L5D3PHI3X1_CM_L3L4_L5D3PHI3X1_wr_en),
.start(VMPROJ_L3L4_L5D3PHI3X1_start),
.done(ME_L3L4_L5D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D3PHI3X2(
.number_in_vmstubin(VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2_number),
.read_add_vmstubin(VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2_read_add),
.vmstubin(VMS_L5D3PHI3X2n5_ME_L3L4_L5D3PHI3X2),
.number_in_vmprojin(VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2_read_add),
.vmprojin(VMPROJ_L3L4_L5D3PHI3X2_ME_L3L4_L5D3PHI3X2),
.matchout(ME_L3L4_L5D3PHI3X2_CM_L3L4_L5D3PHI3X2),
.valid_data(ME_L3L4_L5D3PHI3X2_CM_L3L4_L5D3PHI3X2_wr_en),
.start(VMPROJ_L3L4_L5D3PHI3X2_start),
.done(ME_L3L4_L5D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D4PHI1X1(
.number_in_vmstubin(VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1_number),
.read_add_vmstubin(VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1_read_add),
.vmstubin(VMS_L5D4PHI1X1n5_ME_L3L4_L5D4PHI1X1),
.number_in_vmprojin(VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI1X1_ME_L3L4_L5D4PHI1X1),
.matchout(ME_L3L4_L5D4PHI1X1_CM_L3L4_L5D4PHI1X1),
.valid_data(ME_L3L4_L5D4PHI1X1_CM_L3L4_L5D4PHI1X1_wr_en),
.start(VMPROJ_L3L4_L5D4PHI1X1_start),
.done(ME_L3L4_L5D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D4PHI1X2(
.number_in_vmstubin(VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2_number),
.read_add_vmstubin(VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2_read_add),
.vmstubin(VMS_L5D4PHI1X2n3_ME_L3L4_L5D4PHI1X2),
.number_in_vmprojin(VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI1X2_ME_L3L4_L5D4PHI1X2),
.matchout(ME_L3L4_L5D4PHI1X2_CM_L3L4_L5D4PHI1X2),
.valid_data(ME_L3L4_L5D4PHI1X2_CM_L3L4_L5D4PHI1X2_wr_en),
.start(VMPROJ_L3L4_L5D4PHI1X2_start),
.done(ME_L3L4_L5D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D4PHI2X1(
.number_in_vmstubin(VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1_number),
.read_add_vmstubin(VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1_read_add),
.vmstubin(VMS_L5D4PHI2X1n5_ME_L3L4_L5D4PHI2X1),
.number_in_vmprojin(VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI2X1_ME_L3L4_L5D4PHI2X1),
.matchout(ME_L3L4_L5D4PHI2X1_CM_L3L4_L5D4PHI2X1),
.valid_data(ME_L3L4_L5D4PHI2X1_CM_L3L4_L5D4PHI2X1_wr_en),
.start(VMPROJ_L3L4_L5D4PHI2X1_start),
.done(ME_L3L4_L5D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D4PHI2X2(
.number_in_vmstubin(VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2_number),
.read_add_vmstubin(VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2_read_add),
.vmstubin(VMS_L5D4PHI2X2n3_ME_L3L4_L5D4PHI2X2),
.number_in_vmprojin(VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI2X2_ME_L3L4_L5D4PHI2X2),
.matchout(ME_L3L4_L5D4PHI2X2_CM_L3L4_L5D4PHI2X2),
.valid_data(ME_L3L4_L5D4PHI2X2_CM_L3L4_L5D4PHI2X2_wr_en),
.start(VMPROJ_L3L4_L5D4PHI2X2_start),
.done(ME_L3L4_L5D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D4PHI3X1(
.number_in_vmstubin(VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1_number),
.read_add_vmstubin(VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1_read_add),
.vmstubin(VMS_L5D4PHI3X1n5_ME_L3L4_L5D4PHI3X1),
.number_in_vmprojin(VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI3X1_ME_L3L4_L5D4PHI3X1),
.matchout(ME_L3L4_L5D4PHI3X1_CM_L3L4_L5D4PHI3X1),
.valid_data(ME_L3L4_L5D4PHI3X1_CM_L3L4_L5D4PHI3X1_wr_en),
.start(VMPROJ_L3L4_L5D4PHI3X1_start),
.done(ME_L3L4_L5D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L5D4PHI3X2(
.number_in_vmstubin(VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2_number),
.read_add_vmstubin(VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2_read_add),
.vmstubin(VMS_L5D4PHI3X2n3_ME_L3L4_L5D4PHI3X2),
.number_in_vmprojin(VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2_read_add),
.vmprojin(VMPROJ_L3L4_L5D4PHI3X2_ME_L3L4_L5D4PHI3X2),
.matchout(ME_L3L4_L5D4PHI3X2_CM_L3L4_L5D4PHI3X2),
.valid_data(ME_L3L4_L5D4PHI3X2_CM_L3L4_L5D4PHI3X2_wr_en),
.start(VMPROJ_L3L4_L5D4PHI3X2_start),
.done(ME_L3L4_L5D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D3PHI1X1(
.number_in_vmstubin(VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1_number),
.read_add_vmstubin(VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1_read_add),
.vmstubin(VMS_L6D3PHI1X1n2_ME_L3L4_L6D3PHI1X1),
.number_in_vmprojin(VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI1X1_ME_L3L4_L6D3PHI1X1),
.matchout(ME_L3L4_L6D3PHI1X1_CM_L3L4_L6D3PHI1X1),
.valid_data(ME_L3L4_L6D3PHI1X1_CM_L3L4_L6D3PHI1X1_wr_en),
.start(VMPROJ_L3L4_L6D3PHI1X1_start),
.done(ME_L3L4_L6D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D3PHI1X2(
.number_in_vmstubin(VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2_number),
.read_add_vmstubin(VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2_read_add),
.vmstubin(VMS_L6D3PHI1X2n3_ME_L3L4_L6D3PHI1X2),
.number_in_vmprojin(VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI1X2_ME_L3L4_L6D3PHI1X2),
.matchout(ME_L3L4_L6D3PHI1X2_CM_L3L4_L6D3PHI1X2),
.valid_data(ME_L3L4_L6D3PHI1X2_CM_L3L4_L6D3PHI1X2_wr_en),
.start(VMPROJ_L3L4_L6D3PHI1X2_start),
.done(ME_L3L4_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D3PHI2X1(
.number_in_vmstubin(VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1_number),
.read_add_vmstubin(VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1_read_add),
.vmstubin(VMS_L6D3PHI2X1n3_ME_L3L4_L6D3PHI2X1),
.number_in_vmprojin(VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI2X1_ME_L3L4_L6D3PHI2X1),
.matchout(ME_L3L4_L6D3PHI2X1_CM_L3L4_L6D3PHI2X1),
.valid_data(ME_L3L4_L6D3PHI2X1_CM_L3L4_L6D3PHI2X1_wr_en),
.start(VMPROJ_L3L4_L6D3PHI2X1_start),
.done(ME_L3L4_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D3PHI2X2(
.number_in_vmstubin(VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2_number),
.read_add_vmstubin(VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2_read_add),
.vmstubin(VMS_L6D3PHI2X2n5_ME_L3L4_L6D3PHI2X2),
.number_in_vmprojin(VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI2X2_ME_L3L4_L6D3PHI2X2),
.matchout(ME_L3L4_L6D3PHI2X2_CM_L3L4_L6D3PHI2X2),
.valid_data(ME_L3L4_L6D3PHI2X2_CM_L3L4_L6D3PHI2X2_wr_en),
.start(VMPROJ_L3L4_L6D3PHI2X2_start),
.done(ME_L3L4_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D3PHI3X1(
.number_in_vmstubin(VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1_number),
.read_add_vmstubin(VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1_read_add),
.vmstubin(VMS_L6D3PHI3X1n3_ME_L3L4_L6D3PHI3X1),
.number_in_vmprojin(VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI3X1_ME_L3L4_L6D3PHI3X1),
.matchout(ME_L3L4_L6D3PHI3X1_CM_L3L4_L6D3PHI3X1),
.valid_data(ME_L3L4_L6D3PHI3X1_CM_L3L4_L6D3PHI3X1_wr_en),
.start(VMPROJ_L3L4_L6D3PHI3X1_start),
.done(ME_L3L4_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D3PHI3X2(
.number_in_vmstubin(VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2_number),
.read_add_vmstubin(VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2_read_add),
.vmstubin(VMS_L6D3PHI3X2n5_ME_L3L4_L6D3PHI3X2),
.number_in_vmprojin(VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI3X2_ME_L3L4_L6D3PHI3X2),
.matchout(ME_L3L4_L6D3PHI3X2_CM_L3L4_L6D3PHI3X2),
.valid_data(ME_L3L4_L6D3PHI3X2_CM_L3L4_L6D3PHI3X2_wr_en),
.start(VMPROJ_L3L4_L6D3PHI3X2_start),
.done(ME_L3L4_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D3PHI4X1(
.number_in_vmstubin(VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1_number),
.read_add_vmstubin(VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1_read_add),
.vmstubin(VMS_L6D3PHI4X1n2_ME_L3L4_L6D3PHI4X1),
.number_in_vmprojin(VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI4X1_ME_L3L4_L6D3PHI4X1),
.matchout(ME_L3L4_L6D3PHI4X1_CM_L3L4_L6D3PHI4X1),
.valid_data(ME_L3L4_L6D3PHI4X1_CM_L3L4_L6D3PHI4X1_wr_en),
.start(VMPROJ_L3L4_L6D3PHI4X1_start),
.done(ME_L3L4_L6D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D3PHI4X2(
.number_in_vmstubin(VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2_number),
.read_add_vmstubin(VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2_read_add),
.vmstubin(VMS_L6D3PHI4X2n3_ME_L3L4_L6D3PHI4X2),
.number_in_vmprojin(VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2_read_add),
.vmprojin(VMPROJ_L3L4_L6D3PHI4X2_ME_L3L4_L6D3PHI4X2),
.matchout(ME_L3L4_L6D3PHI4X2_CM_L3L4_L6D3PHI4X2),
.valid_data(ME_L3L4_L6D3PHI4X2_CM_L3L4_L6D3PHI4X2_wr_en),
.start(VMPROJ_L3L4_L6D3PHI4X2_start),
.done(ME_L3L4_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D4PHI1X1(
.number_in_vmstubin(VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1_number),
.read_add_vmstubin(VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1_read_add),
.vmstubin(VMS_L6D4PHI1X1n3_ME_L3L4_L6D4PHI1X1),
.number_in_vmprojin(VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI1X1_ME_L3L4_L6D4PHI1X1),
.matchout(ME_L3L4_L6D4PHI1X1_CM_L3L4_L6D4PHI1X1),
.valid_data(ME_L3L4_L6D4PHI1X1_CM_L3L4_L6D4PHI1X1_wr_en),
.start(VMPROJ_L3L4_L6D4PHI1X1_start),
.done(ME_L3L4_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D4PHI1X2(
.number_in_vmstubin(VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2_number),
.read_add_vmstubin(VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2_read_add),
.vmstubin(VMS_L6D4PHI1X2n3_ME_L3L4_L6D4PHI1X2),
.number_in_vmprojin(VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI1X2_ME_L3L4_L6D4PHI1X2),
.matchout(ME_L3L4_L6D4PHI1X2_CM_L3L4_L6D4PHI1X2),
.valid_data(ME_L3L4_L6D4PHI1X2_CM_L3L4_L6D4PHI1X2_wr_en),
.start(VMPROJ_L3L4_L6D4PHI1X2_start),
.done(ME_L3L4_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D4PHI2X1(
.number_in_vmstubin(VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1_number),
.read_add_vmstubin(VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1_read_add),
.vmstubin(VMS_L6D4PHI2X1n5_ME_L3L4_L6D4PHI2X1),
.number_in_vmprojin(VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI2X1_ME_L3L4_L6D4PHI2X1),
.matchout(ME_L3L4_L6D4PHI2X1_CM_L3L4_L6D4PHI2X1),
.valid_data(ME_L3L4_L6D4PHI2X1_CM_L3L4_L6D4PHI2X1_wr_en),
.start(VMPROJ_L3L4_L6D4PHI2X1_start),
.done(ME_L3L4_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D4PHI2X2(
.number_in_vmstubin(VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2_number),
.read_add_vmstubin(VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2_read_add),
.vmstubin(VMS_L6D4PHI2X2n5_ME_L3L4_L6D4PHI2X2),
.number_in_vmprojin(VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI2X2_ME_L3L4_L6D4PHI2X2),
.matchout(ME_L3L4_L6D4PHI2X2_CM_L3L4_L6D4PHI2X2),
.valid_data(ME_L3L4_L6D4PHI2X2_CM_L3L4_L6D4PHI2X2_wr_en),
.start(VMPROJ_L3L4_L6D4PHI2X2_start),
.done(ME_L3L4_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D4PHI3X1(
.number_in_vmstubin(VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1_number),
.read_add_vmstubin(VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1_read_add),
.vmstubin(VMS_L6D4PHI3X1n5_ME_L3L4_L6D4PHI3X1),
.number_in_vmprojin(VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI3X1_ME_L3L4_L6D4PHI3X1),
.matchout(ME_L3L4_L6D4PHI3X1_CM_L3L4_L6D4PHI3X1),
.valid_data(ME_L3L4_L6D4PHI3X1_CM_L3L4_L6D4PHI3X1_wr_en),
.start(VMPROJ_L3L4_L6D4PHI3X1_start),
.done(ME_L3L4_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D4PHI3X2(
.number_in_vmstubin(VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2_number),
.read_add_vmstubin(VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2_read_add),
.vmstubin(VMS_L6D4PHI3X2n5_ME_L3L4_L6D4PHI3X2),
.number_in_vmprojin(VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI3X2_ME_L3L4_L6D4PHI3X2),
.matchout(ME_L3L4_L6D4PHI3X2_CM_L3L4_L6D4PHI3X2),
.valid_data(ME_L3L4_L6D4PHI3X2_CM_L3L4_L6D4PHI3X2_wr_en),
.start(VMPROJ_L3L4_L6D4PHI3X2_start),
.done(ME_L3L4_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D4PHI4X1(
.number_in_vmstubin(VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1_number),
.read_add_vmstubin(VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1_read_add),
.vmstubin(VMS_L6D4PHI4X1n3_ME_L3L4_L6D4PHI4X1),
.number_in_vmprojin(VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI4X1_ME_L3L4_L6D4PHI4X1),
.matchout(ME_L3L4_L6D4PHI4X1_CM_L3L4_L6D4PHI4X1),
.valid_data(ME_L3L4_L6D4PHI4X1_CM_L3L4_L6D4PHI4X1_wr_en),
.start(VMPROJ_L3L4_L6D4PHI4X1_start),
.done(ME_L3L4_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L3L4_L6D4PHI4X2(
.number_in_vmstubin(VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2_number),
.read_add_vmstubin(VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2_read_add),
.vmstubin(VMS_L6D4PHI4X2n3_ME_L3L4_L6D4PHI4X2),
.number_in_vmprojin(VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2_number),
.read_add_vmprojin(VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2_read_add),
.vmprojin(VMPROJ_L3L4_L6D4PHI4X2_ME_L3L4_L6D4PHI4X2),
.matchout(ME_L3L4_L6D4PHI4X2_CM_L3L4_L6D4PHI4X2),
.valid_data(ME_L3L4_L6D4PHI4X2_CM_L3L4_L6D4PHI4X2_wr_en),
.start(VMPROJ_L3L4_L6D4PHI4X2_start),
.done(ME_L3L4_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D3PHI1X1(
.number_in_vmstubin(VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1_number),
.read_add_vmstubin(VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1_read_add),
.vmstubin(VMS_L3D3PHI1X1n5_ME_L1L2_L3D3PHI1X1),
.number_in_vmprojin(VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI1X1_ME_L1L2_L3D3PHI1X1),
.matchout(ME_L1L2_L3D3PHI1X1_CM_L1L2_L3D3PHI1X1),
.valid_data(ME_L1L2_L3D3PHI1X1_CM_L1L2_L3D3PHI1X1_wr_en),
.start(VMPROJ_L1L2_L3D3PHI1X1_start),
.done(ME_L1L2_L3D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D3PHI1X2(
.number_in_vmstubin(VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2_number),
.read_add_vmstubin(VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2_read_add),
.vmstubin(VMS_L3D3PHI1X2n5_ME_L1L2_L3D3PHI1X2),
.number_in_vmprojin(VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI1X2_ME_L1L2_L3D3PHI1X2),
.matchout(ME_L1L2_L3D3PHI1X2_CM_L1L2_L3D3PHI1X2),
.valid_data(ME_L1L2_L3D3PHI1X2_CM_L1L2_L3D3PHI1X2_wr_en),
.start(VMPROJ_L1L2_L3D3PHI1X2_start),
.done(ME_L1L2_L3D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D3PHI2X1(
.number_in_vmstubin(VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1_number),
.read_add_vmstubin(VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1_read_add),
.vmstubin(VMS_L3D3PHI2X1n5_ME_L1L2_L3D3PHI2X1),
.number_in_vmprojin(VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI2X1_ME_L1L2_L3D3PHI2X1),
.matchout(ME_L1L2_L3D3PHI2X1_CM_L1L2_L3D3PHI2X1),
.valid_data(ME_L1L2_L3D3PHI2X1_CM_L1L2_L3D3PHI2X1_wr_en),
.start(VMPROJ_L1L2_L3D3PHI2X1_start),
.done(ME_L1L2_L3D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D3PHI2X2(
.number_in_vmstubin(VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2_number),
.read_add_vmstubin(VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2_read_add),
.vmstubin(VMS_L3D3PHI2X2n5_ME_L1L2_L3D3PHI2X2),
.number_in_vmprojin(VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI2X2_ME_L1L2_L3D3PHI2X2),
.matchout(ME_L1L2_L3D3PHI2X2_CM_L1L2_L3D3PHI2X2),
.valid_data(ME_L1L2_L3D3PHI2X2_CM_L1L2_L3D3PHI2X2_wr_en),
.start(VMPROJ_L1L2_L3D3PHI2X2_start),
.done(ME_L1L2_L3D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D3PHI3X1(
.number_in_vmstubin(VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1_number),
.read_add_vmstubin(VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1_read_add),
.vmstubin(VMS_L3D3PHI3X1n5_ME_L1L2_L3D3PHI3X1),
.number_in_vmprojin(VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI3X1_ME_L1L2_L3D3PHI3X1),
.matchout(ME_L1L2_L3D3PHI3X1_CM_L1L2_L3D3PHI3X1),
.valid_data(ME_L1L2_L3D3PHI3X1_CM_L1L2_L3D3PHI3X1_wr_en),
.start(VMPROJ_L1L2_L3D3PHI3X1_start),
.done(ME_L1L2_L3D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D3PHI3X2(
.number_in_vmstubin(VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2_number),
.read_add_vmstubin(VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2_read_add),
.vmstubin(VMS_L3D3PHI3X2n5_ME_L1L2_L3D3PHI3X2),
.number_in_vmprojin(VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2_read_add),
.vmprojin(VMPROJ_L1L2_L3D3PHI3X2_ME_L1L2_L3D3PHI3X2),
.matchout(ME_L1L2_L3D3PHI3X2_CM_L1L2_L3D3PHI3X2),
.valid_data(ME_L1L2_L3D3PHI3X2_CM_L1L2_L3D3PHI3X2_wr_en),
.start(VMPROJ_L1L2_L3D3PHI3X2_start),
.done(ME_L1L2_L3D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D4PHI1X1(
.number_in_vmstubin(VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1_number),
.read_add_vmstubin(VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1_read_add),
.vmstubin(VMS_L3D4PHI1X1n5_ME_L1L2_L3D4PHI1X1),
.number_in_vmprojin(VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI1X1_ME_L1L2_L3D4PHI1X1),
.matchout(ME_L1L2_L3D4PHI1X1_CM_L1L2_L3D4PHI1X1),
.valid_data(ME_L1L2_L3D4PHI1X1_CM_L1L2_L3D4PHI1X1_wr_en),
.start(VMPROJ_L1L2_L3D4PHI1X1_start),
.done(ME_L1L2_L3D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D4PHI1X2(
.number_in_vmstubin(VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2_number),
.read_add_vmstubin(VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2_read_add),
.vmstubin(VMS_L3D4PHI1X2n3_ME_L1L2_L3D4PHI1X2),
.number_in_vmprojin(VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI1X2_ME_L1L2_L3D4PHI1X2),
.matchout(ME_L1L2_L3D4PHI1X2_CM_L1L2_L3D4PHI1X2),
.valid_data(ME_L1L2_L3D4PHI1X2_CM_L1L2_L3D4PHI1X2_wr_en),
.start(VMPROJ_L1L2_L3D4PHI1X2_start),
.done(ME_L1L2_L3D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D4PHI2X1(
.number_in_vmstubin(VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1_number),
.read_add_vmstubin(VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1_read_add),
.vmstubin(VMS_L3D4PHI2X1n5_ME_L1L2_L3D4PHI2X1),
.number_in_vmprojin(VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI2X1_ME_L1L2_L3D4PHI2X1),
.matchout(ME_L1L2_L3D4PHI2X1_CM_L1L2_L3D4PHI2X1),
.valid_data(ME_L1L2_L3D4PHI2X1_CM_L1L2_L3D4PHI2X1_wr_en),
.start(VMPROJ_L1L2_L3D4PHI2X1_start),
.done(ME_L1L2_L3D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D4PHI2X2(
.number_in_vmstubin(VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2_number),
.read_add_vmstubin(VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2_read_add),
.vmstubin(VMS_L3D4PHI2X2n3_ME_L1L2_L3D4PHI2X2),
.number_in_vmprojin(VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI2X2_ME_L1L2_L3D4PHI2X2),
.matchout(ME_L1L2_L3D4PHI2X2_CM_L1L2_L3D4PHI2X2),
.valid_data(ME_L1L2_L3D4PHI2X2_CM_L1L2_L3D4PHI2X2_wr_en),
.start(VMPROJ_L1L2_L3D4PHI2X2_start),
.done(ME_L1L2_L3D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D4PHI3X1(
.number_in_vmstubin(VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1_number),
.read_add_vmstubin(VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1_read_add),
.vmstubin(VMS_L3D4PHI3X1n5_ME_L1L2_L3D4PHI3X1),
.number_in_vmprojin(VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI3X1_ME_L1L2_L3D4PHI3X1),
.matchout(ME_L1L2_L3D4PHI3X1_CM_L1L2_L3D4PHI3X1),
.valid_data(ME_L1L2_L3D4PHI3X1_CM_L1L2_L3D4PHI3X1_wr_en),
.start(VMPROJ_L1L2_L3D4PHI3X1_start),
.done(ME_L1L2_L3D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L3D4PHI3X2(
.number_in_vmstubin(VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2_number),
.read_add_vmstubin(VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2_read_add),
.vmstubin(VMS_L3D4PHI3X2n3_ME_L1L2_L3D4PHI3X2),
.number_in_vmprojin(VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2_read_add),
.vmprojin(VMPROJ_L1L2_L3D4PHI3X2_ME_L1L2_L3D4PHI3X2),
.matchout(ME_L1L2_L3D4PHI3X2_CM_L1L2_L3D4PHI3X2),
.valid_data(ME_L1L2_L3D4PHI3X2_CM_L1L2_L3D4PHI3X2_wr_en),
.start(VMPROJ_L1L2_L3D4PHI3X2_start),
.done(ME_L1L2_L3D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D3PHI1X1(
.number_in_vmstubin(VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1_number),
.read_add_vmstubin(VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1_read_add),
.vmstubin(VMS_L4D3PHI1X1n2_ME_L1L2_L4D3PHI1X1),
.number_in_vmprojin(VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI1X1_ME_L1L2_L4D3PHI1X1),
.matchout(ME_L1L2_L4D3PHI1X1_CM_L1L2_L4D3PHI1X1),
.valid_data(ME_L1L2_L4D3PHI1X1_CM_L1L2_L4D3PHI1X1_wr_en),
.start(VMPROJ_L1L2_L4D3PHI1X1_start),
.done(ME_L1L2_L4D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D3PHI1X2(
.number_in_vmstubin(VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2_number),
.read_add_vmstubin(VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2_read_add),
.vmstubin(VMS_L4D3PHI1X2n3_ME_L1L2_L4D3PHI1X2),
.number_in_vmprojin(VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI1X2_ME_L1L2_L4D3PHI1X2),
.matchout(ME_L1L2_L4D3PHI1X2_CM_L1L2_L4D3PHI1X2),
.valid_data(ME_L1L2_L4D3PHI1X2_CM_L1L2_L4D3PHI1X2_wr_en),
.start(VMPROJ_L1L2_L4D3PHI1X2_start),
.done(ME_L1L2_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D3PHI2X1(
.number_in_vmstubin(VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1_number),
.read_add_vmstubin(VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1_read_add),
.vmstubin(VMS_L4D3PHI2X1n3_ME_L1L2_L4D3PHI2X1),
.number_in_vmprojin(VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI2X1_ME_L1L2_L4D3PHI2X1),
.matchout(ME_L1L2_L4D3PHI2X1_CM_L1L2_L4D3PHI2X1),
.valid_data(ME_L1L2_L4D3PHI2X1_CM_L1L2_L4D3PHI2X1_wr_en),
.start(VMPROJ_L1L2_L4D3PHI2X1_start),
.done(ME_L1L2_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D3PHI2X2(
.number_in_vmstubin(VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2_number),
.read_add_vmstubin(VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2_read_add),
.vmstubin(VMS_L4D3PHI2X2n5_ME_L1L2_L4D3PHI2X2),
.number_in_vmprojin(VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI2X2_ME_L1L2_L4D3PHI2X2),
.matchout(ME_L1L2_L4D3PHI2X2_CM_L1L2_L4D3PHI2X2),
.valid_data(ME_L1L2_L4D3PHI2X2_CM_L1L2_L4D3PHI2X2_wr_en),
.start(VMPROJ_L1L2_L4D3PHI2X2_start),
.done(ME_L1L2_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D3PHI3X1(
.number_in_vmstubin(VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1_number),
.read_add_vmstubin(VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1_read_add),
.vmstubin(VMS_L4D3PHI3X1n3_ME_L1L2_L4D3PHI3X1),
.number_in_vmprojin(VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI3X1_ME_L1L2_L4D3PHI3X1),
.matchout(ME_L1L2_L4D3PHI3X1_CM_L1L2_L4D3PHI3X1),
.valid_data(ME_L1L2_L4D3PHI3X1_CM_L1L2_L4D3PHI3X1_wr_en),
.start(VMPROJ_L1L2_L4D3PHI3X1_start),
.done(ME_L1L2_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D3PHI3X2(
.number_in_vmstubin(VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2_number),
.read_add_vmstubin(VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2_read_add),
.vmstubin(VMS_L4D3PHI3X2n5_ME_L1L2_L4D3PHI3X2),
.number_in_vmprojin(VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI3X2_ME_L1L2_L4D3PHI3X2),
.matchout(ME_L1L2_L4D3PHI3X2_CM_L1L2_L4D3PHI3X2),
.valid_data(ME_L1L2_L4D3PHI3X2_CM_L1L2_L4D3PHI3X2_wr_en),
.start(VMPROJ_L1L2_L4D3PHI3X2_start),
.done(ME_L1L2_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D3PHI4X1(
.number_in_vmstubin(VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1_number),
.read_add_vmstubin(VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1_read_add),
.vmstubin(VMS_L4D3PHI4X1n2_ME_L1L2_L4D3PHI4X1),
.number_in_vmprojin(VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI4X1_ME_L1L2_L4D3PHI4X1),
.matchout(ME_L1L2_L4D3PHI4X1_CM_L1L2_L4D3PHI4X1),
.valid_data(ME_L1L2_L4D3PHI4X1_CM_L1L2_L4D3PHI4X1_wr_en),
.start(VMPROJ_L1L2_L4D3PHI4X1_start),
.done(ME_L1L2_L4D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D3PHI4X2(
.number_in_vmstubin(VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2_number),
.read_add_vmstubin(VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2_read_add),
.vmstubin(VMS_L4D3PHI4X2n3_ME_L1L2_L4D3PHI4X2),
.number_in_vmprojin(VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2_read_add),
.vmprojin(VMPROJ_L1L2_L4D3PHI4X2_ME_L1L2_L4D3PHI4X2),
.matchout(ME_L1L2_L4D3PHI4X2_CM_L1L2_L4D3PHI4X2),
.valid_data(ME_L1L2_L4D3PHI4X2_CM_L1L2_L4D3PHI4X2_wr_en),
.start(VMPROJ_L1L2_L4D3PHI4X2_start),
.done(ME_L1L2_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D4PHI1X1(
.number_in_vmstubin(VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1_number),
.read_add_vmstubin(VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1_read_add),
.vmstubin(VMS_L4D4PHI1X1n3_ME_L1L2_L4D4PHI1X1),
.number_in_vmprojin(VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI1X1_ME_L1L2_L4D4PHI1X1),
.matchout(ME_L1L2_L4D4PHI1X1_CM_L1L2_L4D4PHI1X1),
.valid_data(ME_L1L2_L4D4PHI1X1_CM_L1L2_L4D4PHI1X1_wr_en),
.start(VMPROJ_L1L2_L4D4PHI1X1_start),
.done(ME_L1L2_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D4PHI1X2(
.number_in_vmstubin(VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2_number),
.read_add_vmstubin(VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2_read_add),
.vmstubin(VMS_L4D4PHI1X2n3_ME_L1L2_L4D4PHI1X2),
.number_in_vmprojin(VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI1X2_ME_L1L2_L4D4PHI1X2),
.matchout(ME_L1L2_L4D4PHI1X2_CM_L1L2_L4D4PHI1X2),
.valid_data(ME_L1L2_L4D4PHI1X2_CM_L1L2_L4D4PHI1X2_wr_en),
.start(VMPROJ_L1L2_L4D4PHI1X2_start),
.done(ME_L1L2_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D4PHI2X1(
.number_in_vmstubin(VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1_number),
.read_add_vmstubin(VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1_read_add),
.vmstubin(VMS_L4D4PHI2X1n5_ME_L1L2_L4D4PHI2X1),
.number_in_vmprojin(VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI2X1_ME_L1L2_L4D4PHI2X1),
.matchout(ME_L1L2_L4D4PHI2X1_CM_L1L2_L4D4PHI2X1),
.valid_data(ME_L1L2_L4D4PHI2X1_CM_L1L2_L4D4PHI2X1_wr_en),
.start(VMPROJ_L1L2_L4D4PHI2X1_start),
.done(ME_L1L2_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D4PHI2X2(
.number_in_vmstubin(VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2_number),
.read_add_vmstubin(VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2_read_add),
.vmstubin(VMS_L4D4PHI2X2n5_ME_L1L2_L4D4PHI2X2),
.number_in_vmprojin(VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI2X2_ME_L1L2_L4D4PHI2X2),
.matchout(ME_L1L2_L4D4PHI2X2_CM_L1L2_L4D4PHI2X2),
.valid_data(ME_L1L2_L4D4PHI2X2_CM_L1L2_L4D4PHI2X2_wr_en),
.start(VMPROJ_L1L2_L4D4PHI2X2_start),
.done(ME_L1L2_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D4PHI3X1(
.number_in_vmstubin(VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1_number),
.read_add_vmstubin(VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1_read_add),
.vmstubin(VMS_L4D4PHI3X1n5_ME_L1L2_L4D4PHI3X1),
.number_in_vmprojin(VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI3X1_ME_L1L2_L4D4PHI3X1),
.matchout(ME_L1L2_L4D4PHI3X1_CM_L1L2_L4D4PHI3X1),
.valid_data(ME_L1L2_L4D4PHI3X1_CM_L1L2_L4D4PHI3X1_wr_en),
.start(VMPROJ_L1L2_L4D4PHI3X1_start),
.done(ME_L1L2_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D4PHI3X2(
.number_in_vmstubin(VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2_number),
.read_add_vmstubin(VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2_read_add),
.vmstubin(VMS_L4D4PHI3X2n5_ME_L1L2_L4D4PHI3X2),
.number_in_vmprojin(VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI3X2_ME_L1L2_L4D4PHI3X2),
.matchout(ME_L1L2_L4D4PHI3X2_CM_L1L2_L4D4PHI3X2),
.valid_data(ME_L1L2_L4D4PHI3X2_CM_L1L2_L4D4PHI3X2_wr_en),
.start(VMPROJ_L1L2_L4D4PHI3X2_start),
.done(ME_L1L2_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D4PHI4X1(
.number_in_vmstubin(VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1_number),
.read_add_vmstubin(VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1_read_add),
.vmstubin(VMS_L4D4PHI4X1n3_ME_L1L2_L4D4PHI4X1),
.number_in_vmprojin(VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI4X1_ME_L1L2_L4D4PHI4X1),
.matchout(ME_L1L2_L4D4PHI4X1_CM_L1L2_L4D4PHI4X1),
.valid_data(ME_L1L2_L4D4PHI4X1_CM_L1L2_L4D4PHI4X1_wr_en),
.start(VMPROJ_L1L2_L4D4PHI4X1_start),
.done(ME_L1L2_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L4D4PHI4X2(
.number_in_vmstubin(VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2_number),
.read_add_vmstubin(VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2_read_add),
.vmstubin(VMS_L4D4PHI4X2n3_ME_L1L2_L4D4PHI4X2),
.number_in_vmprojin(VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2_read_add),
.vmprojin(VMPROJ_L1L2_L4D4PHI4X2_ME_L1L2_L4D4PHI4X2),
.matchout(ME_L1L2_L4D4PHI4X2_CM_L1L2_L4D4PHI4X2),
.valid_data(ME_L1L2_L4D4PHI4X2_CM_L1L2_L4D4PHI4X2_wr_en),
.start(VMPROJ_L1L2_L4D4PHI4X2_start),
.done(ME_L1L2_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D3PHI1X1(
.number_in_vmstubin(VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1_number),
.read_add_vmstubin(VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1_read_add),
.vmstubin(VMS_L5D3PHI1X1n6_ME_L1L2_L5D3PHI1X1),
.number_in_vmprojin(VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI1X1_ME_L1L2_L5D3PHI1X1),
.matchout(ME_L1L2_L5D3PHI1X1_CM_L1L2_L5D3PHI1X1),
.valid_data(ME_L1L2_L5D3PHI1X1_CM_L1L2_L5D3PHI1X1_wr_en),
.start(VMPROJ_L1L2_L5D3PHI1X1_start),
.done(ME_L1L2_L5D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D3PHI1X2(
.number_in_vmstubin(VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2_number),
.read_add_vmstubin(VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2_read_add),
.vmstubin(VMS_L5D3PHI1X2n6_ME_L1L2_L5D3PHI1X2),
.number_in_vmprojin(VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI1X2_ME_L1L2_L5D3PHI1X2),
.matchout(ME_L1L2_L5D3PHI1X2_CM_L1L2_L5D3PHI1X2),
.valid_data(ME_L1L2_L5D3PHI1X2_CM_L1L2_L5D3PHI1X2_wr_en),
.start(VMPROJ_L1L2_L5D3PHI1X2_start),
.done(ME_L1L2_L5D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D3PHI2X1(
.number_in_vmstubin(VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1_number),
.read_add_vmstubin(VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1_read_add),
.vmstubin(VMS_L5D3PHI2X1n6_ME_L1L2_L5D3PHI2X1),
.number_in_vmprojin(VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI2X1_ME_L1L2_L5D3PHI2X1),
.matchout(ME_L1L2_L5D3PHI2X1_CM_L1L2_L5D3PHI2X1),
.valid_data(ME_L1L2_L5D3PHI2X1_CM_L1L2_L5D3PHI2X1_wr_en),
.start(VMPROJ_L1L2_L5D3PHI2X1_start),
.done(ME_L1L2_L5D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D3PHI2X2(
.number_in_vmstubin(VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2_number),
.read_add_vmstubin(VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2_read_add),
.vmstubin(VMS_L5D3PHI2X2n6_ME_L1L2_L5D3PHI2X2),
.number_in_vmprojin(VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI2X2_ME_L1L2_L5D3PHI2X2),
.matchout(ME_L1L2_L5D3PHI2X2_CM_L1L2_L5D3PHI2X2),
.valid_data(ME_L1L2_L5D3PHI2X2_CM_L1L2_L5D3PHI2X2_wr_en),
.start(VMPROJ_L1L2_L5D3PHI2X2_start),
.done(ME_L1L2_L5D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D3PHI3X1(
.number_in_vmstubin(VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1_number),
.read_add_vmstubin(VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1_read_add),
.vmstubin(VMS_L5D3PHI3X1n6_ME_L1L2_L5D3PHI3X1),
.number_in_vmprojin(VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI3X1_ME_L1L2_L5D3PHI3X1),
.matchout(ME_L1L2_L5D3PHI3X1_CM_L1L2_L5D3PHI3X1),
.valid_data(ME_L1L2_L5D3PHI3X1_CM_L1L2_L5D3PHI3X1_wr_en),
.start(VMPROJ_L1L2_L5D3PHI3X1_start),
.done(ME_L1L2_L5D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D3PHI3X2(
.number_in_vmstubin(VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2_number),
.read_add_vmstubin(VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2_read_add),
.vmstubin(VMS_L5D3PHI3X2n6_ME_L1L2_L5D3PHI3X2),
.number_in_vmprojin(VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2_read_add),
.vmprojin(VMPROJ_L1L2_L5D3PHI3X2_ME_L1L2_L5D3PHI3X2),
.matchout(ME_L1L2_L5D3PHI3X2_CM_L1L2_L5D3PHI3X2),
.valid_data(ME_L1L2_L5D3PHI3X2_CM_L1L2_L5D3PHI3X2_wr_en),
.start(VMPROJ_L1L2_L5D3PHI3X2_start),
.done(ME_L1L2_L5D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D4PHI1X1(
.number_in_vmstubin(VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1_number),
.read_add_vmstubin(VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1_read_add),
.vmstubin(VMS_L5D4PHI1X1n6_ME_L1L2_L5D4PHI1X1),
.number_in_vmprojin(VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI1X1_ME_L1L2_L5D4PHI1X1),
.matchout(ME_L1L2_L5D4PHI1X1_CM_L1L2_L5D4PHI1X1),
.valid_data(ME_L1L2_L5D4PHI1X1_CM_L1L2_L5D4PHI1X1_wr_en),
.start(VMPROJ_L1L2_L5D4PHI1X1_start),
.done(ME_L1L2_L5D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D4PHI1X2(
.number_in_vmstubin(VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2_number),
.read_add_vmstubin(VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2_read_add),
.vmstubin(VMS_L5D4PHI1X2n4_ME_L1L2_L5D4PHI1X2),
.number_in_vmprojin(VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI1X2_ME_L1L2_L5D4PHI1X2),
.matchout(ME_L1L2_L5D4PHI1X2_CM_L1L2_L5D4PHI1X2),
.valid_data(ME_L1L2_L5D4PHI1X2_CM_L1L2_L5D4PHI1X2_wr_en),
.start(VMPROJ_L1L2_L5D4PHI1X2_start),
.done(ME_L1L2_L5D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D4PHI2X1(
.number_in_vmstubin(VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1_number),
.read_add_vmstubin(VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1_read_add),
.vmstubin(VMS_L5D4PHI2X1n6_ME_L1L2_L5D4PHI2X1),
.number_in_vmprojin(VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI2X1_ME_L1L2_L5D4PHI2X1),
.matchout(ME_L1L2_L5D4PHI2X1_CM_L1L2_L5D4PHI2X1),
.valid_data(ME_L1L2_L5D4PHI2X1_CM_L1L2_L5D4PHI2X1_wr_en),
.start(VMPROJ_L1L2_L5D4PHI2X1_start),
.done(ME_L1L2_L5D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D4PHI2X2(
.number_in_vmstubin(VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2_number),
.read_add_vmstubin(VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2_read_add),
.vmstubin(VMS_L5D4PHI2X2n4_ME_L1L2_L5D4PHI2X2),
.number_in_vmprojin(VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI2X2_ME_L1L2_L5D4PHI2X2),
.matchout(ME_L1L2_L5D4PHI2X2_CM_L1L2_L5D4PHI2X2),
.valid_data(ME_L1L2_L5D4PHI2X2_CM_L1L2_L5D4PHI2X2_wr_en),
.start(VMPROJ_L1L2_L5D4PHI2X2_start),
.done(ME_L1L2_L5D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D4PHI3X1(
.number_in_vmstubin(VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1_number),
.read_add_vmstubin(VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1_read_add),
.vmstubin(VMS_L5D4PHI3X1n6_ME_L1L2_L5D4PHI3X1),
.number_in_vmprojin(VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI3X1_ME_L1L2_L5D4PHI3X1),
.matchout(ME_L1L2_L5D4PHI3X1_CM_L1L2_L5D4PHI3X1),
.valid_data(ME_L1L2_L5D4PHI3X1_CM_L1L2_L5D4PHI3X1_wr_en),
.start(VMPROJ_L1L2_L5D4PHI3X1_start),
.done(ME_L1L2_L5D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L5D4PHI3X2(
.number_in_vmstubin(VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2_number),
.read_add_vmstubin(VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2_read_add),
.vmstubin(VMS_L5D4PHI3X2n4_ME_L1L2_L5D4PHI3X2),
.number_in_vmprojin(VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2_read_add),
.vmprojin(VMPROJ_L1L2_L5D4PHI3X2_ME_L1L2_L5D4PHI3X2),
.matchout(ME_L1L2_L5D4PHI3X2_CM_L1L2_L5D4PHI3X2),
.valid_data(ME_L1L2_L5D4PHI3X2_CM_L1L2_L5D4PHI3X2_wr_en),
.start(VMPROJ_L1L2_L5D4PHI3X2_start),
.done(ME_L1L2_L5D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D3PHI1X1(
.number_in_vmstubin(VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1_number),
.read_add_vmstubin(VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1_read_add),
.vmstubin(VMS_L6D3PHI1X1n3_ME_L1L2_L6D3PHI1X1),
.number_in_vmprojin(VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI1X1_ME_L1L2_L6D3PHI1X1),
.matchout(ME_L1L2_L6D3PHI1X1_CM_L1L2_L6D3PHI1X1),
.valid_data(ME_L1L2_L6D3PHI1X1_CM_L1L2_L6D3PHI1X1_wr_en),
.start(VMPROJ_L1L2_L6D3PHI1X1_start),
.done(ME_L1L2_L6D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D3PHI1X2(
.number_in_vmstubin(VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2_number),
.read_add_vmstubin(VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2_read_add),
.vmstubin(VMS_L6D3PHI1X2n4_ME_L1L2_L6D3PHI1X2),
.number_in_vmprojin(VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI1X2_ME_L1L2_L6D3PHI1X2),
.matchout(ME_L1L2_L6D3PHI1X2_CM_L1L2_L6D3PHI1X2),
.valid_data(ME_L1L2_L6D3PHI1X2_CM_L1L2_L6D3PHI1X2_wr_en),
.start(VMPROJ_L1L2_L6D3PHI1X2_start),
.done(ME_L1L2_L6D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D3PHI2X1(
.number_in_vmstubin(VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1_number),
.read_add_vmstubin(VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1_read_add),
.vmstubin(VMS_L6D3PHI2X1n4_ME_L1L2_L6D3PHI2X1),
.number_in_vmprojin(VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI2X1_ME_L1L2_L6D3PHI2X1),
.matchout(ME_L1L2_L6D3PHI2X1_CM_L1L2_L6D3PHI2X1),
.valid_data(ME_L1L2_L6D3PHI2X1_CM_L1L2_L6D3PHI2X1_wr_en),
.start(VMPROJ_L1L2_L6D3PHI2X1_start),
.done(ME_L1L2_L6D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D3PHI2X2(
.number_in_vmstubin(VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2_number),
.read_add_vmstubin(VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2_read_add),
.vmstubin(VMS_L6D3PHI2X2n6_ME_L1L2_L6D3PHI2X2),
.number_in_vmprojin(VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI2X2_ME_L1L2_L6D3PHI2X2),
.matchout(ME_L1L2_L6D3PHI2X2_CM_L1L2_L6D3PHI2X2),
.valid_data(ME_L1L2_L6D3PHI2X2_CM_L1L2_L6D3PHI2X2_wr_en),
.start(VMPROJ_L1L2_L6D3PHI2X2_start),
.done(ME_L1L2_L6D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D3PHI3X1(
.number_in_vmstubin(VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1_number),
.read_add_vmstubin(VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1_read_add),
.vmstubin(VMS_L6D3PHI3X1n4_ME_L1L2_L6D3PHI3X1),
.number_in_vmprojin(VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI3X1_ME_L1L2_L6D3PHI3X1),
.matchout(ME_L1L2_L6D3PHI3X1_CM_L1L2_L6D3PHI3X1),
.valid_data(ME_L1L2_L6D3PHI3X1_CM_L1L2_L6D3PHI3X1_wr_en),
.start(VMPROJ_L1L2_L6D3PHI3X1_start),
.done(ME_L1L2_L6D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D3PHI3X2(
.number_in_vmstubin(VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2_number),
.read_add_vmstubin(VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2_read_add),
.vmstubin(VMS_L6D3PHI3X2n6_ME_L1L2_L6D3PHI3X2),
.number_in_vmprojin(VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI3X2_ME_L1L2_L6D3PHI3X2),
.matchout(ME_L1L2_L6D3PHI3X2_CM_L1L2_L6D3PHI3X2),
.valid_data(ME_L1L2_L6D3PHI3X2_CM_L1L2_L6D3PHI3X2_wr_en),
.start(VMPROJ_L1L2_L6D3PHI3X2_start),
.done(ME_L1L2_L6D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D3PHI4X1(
.number_in_vmstubin(VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1_number),
.read_add_vmstubin(VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1_read_add),
.vmstubin(VMS_L6D3PHI4X1n3_ME_L1L2_L6D3PHI4X1),
.number_in_vmprojin(VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI4X1_ME_L1L2_L6D3PHI4X1),
.matchout(ME_L1L2_L6D3PHI4X1_CM_L1L2_L6D3PHI4X1),
.valid_data(ME_L1L2_L6D3PHI4X1_CM_L1L2_L6D3PHI4X1_wr_en),
.start(VMPROJ_L1L2_L6D3PHI4X1_start),
.done(ME_L1L2_L6D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D3PHI4X2(
.number_in_vmstubin(VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2_number),
.read_add_vmstubin(VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2_read_add),
.vmstubin(VMS_L6D3PHI4X2n4_ME_L1L2_L6D3PHI4X2),
.number_in_vmprojin(VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2_read_add),
.vmprojin(VMPROJ_L1L2_L6D3PHI4X2_ME_L1L2_L6D3PHI4X2),
.matchout(ME_L1L2_L6D3PHI4X2_CM_L1L2_L6D3PHI4X2),
.valid_data(ME_L1L2_L6D3PHI4X2_CM_L1L2_L6D3PHI4X2_wr_en),
.start(VMPROJ_L1L2_L6D3PHI4X2_start),
.done(ME_L1L2_L6D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D4PHI1X1(
.number_in_vmstubin(VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1_number),
.read_add_vmstubin(VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1_read_add),
.vmstubin(VMS_L6D4PHI1X1n4_ME_L1L2_L6D4PHI1X1),
.number_in_vmprojin(VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI1X1_ME_L1L2_L6D4PHI1X1),
.matchout(ME_L1L2_L6D4PHI1X1_CM_L1L2_L6D4PHI1X1),
.valid_data(ME_L1L2_L6D4PHI1X1_CM_L1L2_L6D4PHI1X1_wr_en),
.start(VMPROJ_L1L2_L6D4PHI1X1_start),
.done(ME_L1L2_L6D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D4PHI1X2(
.number_in_vmstubin(VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2_number),
.read_add_vmstubin(VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2_read_add),
.vmstubin(VMS_L6D4PHI1X2n4_ME_L1L2_L6D4PHI1X2),
.number_in_vmprojin(VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI1X2_ME_L1L2_L6D4PHI1X2),
.matchout(ME_L1L2_L6D4PHI1X2_CM_L1L2_L6D4PHI1X2),
.valid_data(ME_L1L2_L6D4PHI1X2_CM_L1L2_L6D4PHI1X2_wr_en),
.start(VMPROJ_L1L2_L6D4PHI1X2_start),
.done(ME_L1L2_L6D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D4PHI2X1(
.number_in_vmstubin(VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1_number),
.read_add_vmstubin(VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1_read_add),
.vmstubin(VMS_L6D4PHI2X1n6_ME_L1L2_L6D4PHI2X1),
.number_in_vmprojin(VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI2X1_ME_L1L2_L6D4PHI2X1),
.matchout(ME_L1L2_L6D4PHI2X1_CM_L1L2_L6D4PHI2X1),
.valid_data(ME_L1L2_L6D4PHI2X1_CM_L1L2_L6D4PHI2X1_wr_en),
.start(VMPROJ_L1L2_L6D4PHI2X1_start),
.done(ME_L1L2_L6D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D4PHI2X2(
.number_in_vmstubin(VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2_number),
.read_add_vmstubin(VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2_read_add),
.vmstubin(VMS_L6D4PHI2X2n6_ME_L1L2_L6D4PHI2X2),
.number_in_vmprojin(VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI2X2_ME_L1L2_L6D4PHI2X2),
.matchout(ME_L1L2_L6D4PHI2X2_CM_L1L2_L6D4PHI2X2),
.valid_data(ME_L1L2_L6D4PHI2X2_CM_L1L2_L6D4PHI2X2_wr_en),
.start(VMPROJ_L1L2_L6D4PHI2X2_start),
.done(ME_L1L2_L6D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D4PHI3X1(
.number_in_vmstubin(VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1_number),
.read_add_vmstubin(VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1_read_add),
.vmstubin(VMS_L6D4PHI3X1n6_ME_L1L2_L6D4PHI3X1),
.number_in_vmprojin(VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI3X1_ME_L1L2_L6D4PHI3X1),
.matchout(ME_L1L2_L6D4PHI3X1_CM_L1L2_L6D4PHI3X1),
.valid_data(ME_L1L2_L6D4PHI3X1_CM_L1L2_L6D4PHI3X1_wr_en),
.start(VMPROJ_L1L2_L6D4PHI3X1_start),
.done(ME_L1L2_L6D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D4PHI3X2(
.number_in_vmstubin(VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2_number),
.read_add_vmstubin(VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2_read_add),
.vmstubin(VMS_L6D4PHI3X2n6_ME_L1L2_L6D4PHI3X2),
.number_in_vmprojin(VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI3X2_ME_L1L2_L6D4PHI3X2),
.matchout(ME_L1L2_L6D4PHI3X2_CM_L1L2_L6D4PHI3X2),
.valid_data(ME_L1L2_L6D4PHI3X2_CM_L1L2_L6D4PHI3X2_wr_en),
.start(VMPROJ_L1L2_L6D4PHI3X2_start),
.done(ME_L1L2_L6D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D4PHI4X1(
.number_in_vmstubin(VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1_number),
.read_add_vmstubin(VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1_read_add),
.vmstubin(VMS_L6D4PHI4X1n4_ME_L1L2_L6D4PHI4X1),
.number_in_vmprojin(VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI4X1_ME_L1L2_L6D4PHI4X1),
.matchout(ME_L1L2_L6D4PHI4X1_CM_L1L2_L6D4PHI4X1),
.valid_data(ME_L1L2_L6D4PHI4X1_CM_L1L2_L6D4PHI4X1_wr_en),
.start(VMPROJ_L1L2_L6D4PHI4X1_start),
.done(ME_L1L2_L6D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L1L2_L6D4PHI4X2(
.number_in_vmstubin(VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2_number),
.read_add_vmstubin(VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2_read_add),
.vmstubin(VMS_L6D4PHI4X2n4_ME_L1L2_L6D4PHI4X2),
.number_in_vmprojin(VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2_number),
.read_add_vmprojin(VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2_read_add),
.vmprojin(VMPROJ_L1L2_L6D4PHI4X2_ME_L1L2_L6D4PHI4X2),
.matchout(ME_L1L2_L6D4PHI4X2_CM_L1L2_L6D4PHI4X2),
.valid_data(ME_L1L2_L6D4PHI4X2_CM_L1L2_L6D4PHI4X2_wr_en),
.start(VMPROJ_L1L2_L6D4PHI4X2_start),
.done(ME_L1L2_L6D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D3PHI1X1(
.number_in_vmstubin(VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1_number),
.read_add_vmstubin(VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1_read_add),
.vmstubin(VMS_L1D3PHI1X1n8_ME_L5L6_L1D3PHI1X1),
.number_in_vmprojin(VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI1X1_ME_L5L6_L1D3PHI1X1),
.matchout(ME_L5L6_L1D3PHI1X1_CM_L5L6_L1D3PHI1X1),
.valid_data(ME_L5L6_L1D3PHI1X1_CM_L5L6_L1D3PHI1X1_wr_en),
.start(VMPROJ_L5L6_L1D3PHI1X1_start),
.done(ME_L5L6_L1D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D3PHI1X2(
.number_in_vmstubin(VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2_number),
.read_add_vmstubin(VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2_read_add),
.vmstubin(VMS_L1D3PHI1X2n8_ME_L5L6_L1D3PHI1X2),
.number_in_vmprojin(VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI1X2_ME_L5L6_L1D3PHI1X2),
.matchout(ME_L5L6_L1D3PHI1X2_CM_L5L6_L1D3PHI1X2),
.valid_data(ME_L5L6_L1D3PHI1X2_CM_L5L6_L1D3PHI1X2_wr_en),
.start(VMPROJ_L5L6_L1D3PHI1X2_start),
.done(ME_L5L6_L1D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D3PHI2X1(
.number_in_vmstubin(VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1_number),
.read_add_vmstubin(VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1_read_add),
.vmstubin(VMS_L1D3PHI2X1n8_ME_L5L6_L1D3PHI2X1),
.number_in_vmprojin(VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI2X1_ME_L5L6_L1D3PHI2X1),
.matchout(ME_L5L6_L1D3PHI2X1_CM_L5L6_L1D3PHI2X1),
.valid_data(ME_L5L6_L1D3PHI2X1_CM_L5L6_L1D3PHI2X1_wr_en),
.start(VMPROJ_L5L6_L1D3PHI2X1_start),
.done(ME_L5L6_L1D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D3PHI2X2(
.number_in_vmstubin(VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2_number),
.read_add_vmstubin(VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2_read_add),
.vmstubin(VMS_L1D3PHI2X2n8_ME_L5L6_L1D3PHI2X2),
.number_in_vmprojin(VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI2X2_ME_L5L6_L1D3PHI2X2),
.matchout(ME_L5L6_L1D3PHI2X2_CM_L5L6_L1D3PHI2X2),
.valid_data(ME_L5L6_L1D3PHI2X2_CM_L5L6_L1D3PHI2X2_wr_en),
.start(VMPROJ_L5L6_L1D3PHI2X2_start),
.done(ME_L5L6_L1D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D3PHI3X1(
.number_in_vmstubin(VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1_number),
.read_add_vmstubin(VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1_read_add),
.vmstubin(VMS_L1D3PHI3X1n8_ME_L5L6_L1D3PHI3X1),
.number_in_vmprojin(VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI3X1_ME_L5L6_L1D3PHI3X1),
.matchout(ME_L5L6_L1D3PHI3X1_CM_L5L6_L1D3PHI3X1),
.valid_data(ME_L5L6_L1D3PHI3X1_CM_L5L6_L1D3PHI3X1_wr_en),
.start(VMPROJ_L5L6_L1D3PHI3X1_start),
.done(ME_L5L6_L1D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D3PHI3X2(
.number_in_vmstubin(VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2_number),
.read_add_vmstubin(VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2_read_add),
.vmstubin(VMS_L1D3PHI3X2n8_ME_L5L6_L1D3PHI3X2),
.number_in_vmprojin(VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2_read_add),
.vmprojin(VMPROJ_L5L6_L1D3PHI3X2_ME_L5L6_L1D3PHI3X2),
.matchout(ME_L5L6_L1D3PHI3X2_CM_L5L6_L1D3PHI3X2),
.valid_data(ME_L5L6_L1D3PHI3X2_CM_L5L6_L1D3PHI3X2_wr_en),
.start(VMPROJ_L5L6_L1D3PHI3X2_start),
.done(ME_L5L6_L1D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D4PHI1X1(
.number_in_vmstubin(VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1_number),
.read_add_vmstubin(VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1_read_add),
.vmstubin(VMS_L1D4PHI1X1n4_ME_L5L6_L1D4PHI1X1),
.number_in_vmprojin(VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI1X1_ME_L5L6_L1D4PHI1X1),
.matchout(ME_L5L6_L1D4PHI1X1_CM_L5L6_L1D4PHI1X1),
.valid_data(ME_L5L6_L1D4PHI1X1_CM_L5L6_L1D4PHI1X1_wr_en),
.start(VMPROJ_L5L6_L1D4PHI1X1_start),
.done(ME_L5L6_L1D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D4PHI1X2(
.number_in_vmstubin(VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2_number),
.read_add_vmstubin(VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2_read_add),
.vmstubin(VMS_L1D4PHI1X2n2_ME_L5L6_L1D4PHI1X2),
.number_in_vmprojin(VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI1X2_ME_L5L6_L1D4PHI1X2),
.matchout(ME_L5L6_L1D4PHI1X2_CM_L5L6_L1D4PHI1X2),
.valid_data(ME_L5L6_L1D4PHI1X2_CM_L5L6_L1D4PHI1X2_wr_en),
.start(VMPROJ_L5L6_L1D4PHI1X2_start),
.done(ME_L5L6_L1D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D4PHI2X1(
.number_in_vmstubin(VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1_number),
.read_add_vmstubin(VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1_read_add),
.vmstubin(VMS_L1D4PHI2X1n4_ME_L5L6_L1D4PHI2X1),
.number_in_vmprojin(VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI2X1_ME_L5L6_L1D4PHI2X1),
.matchout(ME_L5L6_L1D4PHI2X1_CM_L5L6_L1D4PHI2X1),
.valid_data(ME_L5L6_L1D4PHI2X1_CM_L5L6_L1D4PHI2X1_wr_en),
.start(VMPROJ_L5L6_L1D4PHI2X1_start),
.done(ME_L5L6_L1D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D4PHI2X2(
.number_in_vmstubin(VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2_number),
.read_add_vmstubin(VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2_read_add),
.vmstubin(VMS_L1D4PHI2X2n2_ME_L5L6_L1D4PHI2X2),
.number_in_vmprojin(VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI2X2_ME_L5L6_L1D4PHI2X2),
.matchout(ME_L5L6_L1D4PHI2X2_CM_L5L6_L1D4PHI2X2),
.valid_data(ME_L5L6_L1D4PHI2X2_CM_L5L6_L1D4PHI2X2_wr_en),
.start(VMPROJ_L5L6_L1D4PHI2X2_start),
.done(ME_L5L6_L1D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D4PHI3X1(
.number_in_vmstubin(VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1_number),
.read_add_vmstubin(VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1_read_add),
.vmstubin(VMS_L1D4PHI3X1n4_ME_L5L6_L1D4PHI3X1),
.number_in_vmprojin(VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI3X1_ME_L5L6_L1D4PHI3X1),
.matchout(ME_L5L6_L1D4PHI3X1_CM_L5L6_L1D4PHI3X1),
.valid_data(ME_L5L6_L1D4PHI3X1_CM_L5L6_L1D4PHI3X1_wr_en),
.start(VMPROJ_L5L6_L1D4PHI3X1_start),
.done(ME_L5L6_L1D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L1D4PHI3X2(
.number_in_vmstubin(VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2_number),
.read_add_vmstubin(VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2_read_add),
.vmstubin(VMS_L1D4PHI3X2n2_ME_L5L6_L1D4PHI3X2),
.number_in_vmprojin(VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2_read_add),
.vmprojin(VMPROJ_L5L6_L1D4PHI3X2_ME_L5L6_L1D4PHI3X2),
.matchout(ME_L5L6_L1D4PHI3X2_CM_L5L6_L1D4PHI3X2),
.valid_data(ME_L5L6_L1D4PHI3X2_CM_L5L6_L1D4PHI3X2_wr_en),
.start(VMPROJ_L5L6_L1D4PHI3X2_start),
.done(ME_L5L6_L1D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D3PHI1X1(
.number_in_vmstubin(VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1_number),
.read_add_vmstubin(VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1_read_add),
.vmstubin(VMS_L2D3PHI1X1n3_ME_L5L6_L2D3PHI1X1),
.number_in_vmprojin(VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI1X1_ME_L5L6_L2D3PHI1X1),
.matchout(ME_L5L6_L2D3PHI1X1_CM_L5L6_L2D3PHI1X1),
.valid_data(ME_L5L6_L2D3PHI1X1_CM_L5L6_L2D3PHI1X1_wr_en),
.start(VMPROJ_L5L6_L2D3PHI1X1_start),
.done(ME_L5L6_L2D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D3PHI1X2(
.number_in_vmstubin(VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2_number),
.read_add_vmstubin(VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2_read_add),
.vmstubin(VMS_L2D3PHI1X2n4_ME_L5L6_L2D3PHI1X2),
.number_in_vmprojin(VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI1X2_ME_L5L6_L2D3PHI1X2),
.matchout(ME_L5L6_L2D3PHI1X2_CM_L5L6_L2D3PHI1X2),
.valid_data(ME_L5L6_L2D3PHI1X2_CM_L5L6_L2D3PHI1X2_wr_en),
.start(VMPROJ_L5L6_L2D3PHI1X2_start),
.done(ME_L5L6_L2D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D3PHI2X1(
.number_in_vmstubin(VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1_number),
.read_add_vmstubin(VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1_read_add),
.vmstubin(VMS_L2D3PHI2X1n4_ME_L5L6_L2D3PHI2X1),
.number_in_vmprojin(VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI2X1_ME_L5L6_L2D3PHI2X1),
.matchout(ME_L5L6_L2D3PHI2X1_CM_L5L6_L2D3PHI2X1),
.valid_data(ME_L5L6_L2D3PHI2X1_CM_L5L6_L2D3PHI2X1_wr_en),
.start(VMPROJ_L5L6_L2D3PHI2X1_start),
.done(ME_L5L6_L2D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D3PHI2X2(
.number_in_vmstubin(VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2_number),
.read_add_vmstubin(VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2_read_add),
.vmstubin(VMS_L2D3PHI2X2n6_ME_L5L6_L2D3PHI2X2),
.number_in_vmprojin(VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI2X2_ME_L5L6_L2D3PHI2X2),
.matchout(ME_L5L6_L2D3PHI2X2_CM_L5L6_L2D3PHI2X2),
.valid_data(ME_L5L6_L2D3PHI2X2_CM_L5L6_L2D3PHI2X2_wr_en),
.start(VMPROJ_L5L6_L2D3PHI2X2_start),
.done(ME_L5L6_L2D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D3PHI3X1(
.number_in_vmstubin(VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1_number),
.read_add_vmstubin(VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1_read_add),
.vmstubin(VMS_L2D3PHI3X1n4_ME_L5L6_L2D3PHI3X1),
.number_in_vmprojin(VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI3X1_ME_L5L6_L2D3PHI3X1),
.matchout(ME_L5L6_L2D3PHI3X1_CM_L5L6_L2D3PHI3X1),
.valid_data(ME_L5L6_L2D3PHI3X1_CM_L5L6_L2D3PHI3X1_wr_en),
.start(VMPROJ_L5L6_L2D3PHI3X1_start),
.done(ME_L5L6_L2D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D3PHI3X2(
.number_in_vmstubin(VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2_number),
.read_add_vmstubin(VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2_read_add),
.vmstubin(VMS_L2D3PHI3X2n6_ME_L5L6_L2D3PHI3X2),
.number_in_vmprojin(VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI3X2_ME_L5L6_L2D3PHI3X2),
.matchout(ME_L5L6_L2D3PHI3X2_CM_L5L6_L2D3PHI3X2),
.valid_data(ME_L5L6_L2D3PHI3X2_CM_L5L6_L2D3PHI3X2_wr_en),
.start(VMPROJ_L5L6_L2D3PHI3X2_start),
.done(ME_L5L6_L2D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D3PHI4X1(
.number_in_vmstubin(VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1_number),
.read_add_vmstubin(VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1_read_add),
.vmstubin(VMS_L2D3PHI4X1n3_ME_L5L6_L2D3PHI4X1),
.number_in_vmprojin(VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI4X1_ME_L5L6_L2D3PHI4X1),
.matchout(ME_L5L6_L2D3PHI4X1_CM_L5L6_L2D3PHI4X1),
.valid_data(ME_L5L6_L2D3PHI4X1_CM_L5L6_L2D3PHI4X1_wr_en),
.start(VMPROJ_L5L6_L2D3PHI4X1_start),
.done(ME_L5L6_L2D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D3PHI4X2(
.number_in_vmstubin(VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2_number),
.read_add_vmstubin(VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2_read_add),
.vmstubin(VMS_L2D3PHI4X2n4_ME_L5L6_L2D3PHI4X2),
.number_in_vmprojin(VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2_read_add),
.vmprojin(VMPROJ_L5L6_L2D3PHI4X2_ME_L5L6_L2D3PHI4X2),
.matchout(ME_L5L6_L2D3PHI4X2_CM_L5L6_L2D3PHI4X2),
.valid_data(ME_L5L6_L2D3PHI4X2_CM_L5L6_L2D3PHI4X2_wr_en),
.start(VMPROJ_L5L6_L2D3PHI4X2_start),
.done(ME_L5L6_L2D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D4PHI1X1(
.number_in_vmstubin(VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1_number),
.read_add_vmstubin(VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1_read_add),
.vmstubin(VMS_L2D4PHI1X1n4_ME_L5L6_L2D4PHI1X1),
.number_in_vmprojin(VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI1X1_ME_L5L6_L2D4PHI1X1),
.matchout(ME_L5L6_L2D4PHI1X1_CM_L5L6_L2D4PHI1X1),
.valid_data(ME_L5L6_L2D4PHI1X1_CM_L5L6_L2D4PHI1X1_wr_en),
.start(VMPROJ_L5L6_L2D4PHI1X1_start),
.done(ME_L5L6_L2D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D4PHI1X2(
.number_in_vmstubin(VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2_number),
.read_add_vmstubin(VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2_read_add),
.vmstubin(VMS_L2D4PHI1X2n4_ME_L5L6_L2D4PHI1X2),
.number_in_vmprojin(VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI1X2_ME_L5L6_L2D4PHI1X2),
.matchout(ME_L5L6_L2D4PHI1X2_CM_L5L6_L2D4PHI1X2),
.valid_data(ME_L5L6_L2D4PHI1X2_CM_L5L6_L2D4PHI1X2_wr_en),
.start(VMPROJ_L5L6_L2D4PHI1X2_start),
.done(ME_L5L6_L2D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D4PHI2X1(
.number_in_vmstubin(VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1_number),
.read_add_vmstubin(VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1_read_add),
.vmstubin(VMS_L2D4PHI2X1n6_ME_L5L6_L2D4PHI2X1),
.number_in_vmprojin(VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI2X1_ME_L5L6_L2D4PHI2X1),
.matchout(ME_L5L6_L2D4PHI2X1_CM_L5L6_L2D4PHI2X1),
.valid_data(ME_L5L6_L2D4PHI2X1_CM_L5L6_L2D4PHI2X1_wr_en),
.start(VMPROJ_L5L6_L2D4PHI2X1_start),
.done(ME_L5L6_L2D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D4PHI2X2(
.number_in_vmstubin(VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2_number),
.read_add_vmstubin(VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2_read_add),
.vmstubin(VMS_L2D4PHI2X2n6_ME_L5L6_L2D4PHI2X2),
.number_in_vmprojin(VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI2X2_ME_L5L6_L2D4PHI2X2),
.matchout(ME_L5L6_L2D4PHI2X2_CM_L5L6_L2D4PHI2X2),
.valid_data(ME_L5L6_L2D4PHI2X2_CM_L5L6_L2D4PHI2X2_wr_en),
.start(VMPROJ_L5L6_L2D4PHI2X2_start),
.done(ME_L5L6_L2D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D4PHI3X1(
.number_in_vmstubin(VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1_number),
.read_add_vmstubin(VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1_read_add),
.vmstubin(VMS_L2D4PHI3X1n6_ME_L5L6_L2D4PHI3X1),
.number_in_vmprojin(VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI3X1_ME_L5L6_L2D4PHI3X1),
.matchout(ME_L5L6_L2D4PHI3X1_CM_L5L6_L2D4PHI3X1),
.valid_data(ME_L5L6_L2D4PHI3X1_CM_L5L6_L2D4PHI3X1_wr_en),
.start(VMPROJ_L5L6_L2D4PHI3X1_start),
.done(ME_L5L6_L2D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D4PHI3X2(
.number_in_vmstubin(VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2_number),
.read_add_vmstubin(VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2_read_add),
.vmstubin(VMS_L2D4PHI3X2n6_ME_L5L6_L2D4PHI3X2),
.number_in_vmprojin(VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI3X2_ME_L5L6_L2D4PHI3X2),
.matchout(ME_L5L6_L2D4PHI3X2_CM_L5L6_L2D4PHI3X2),
.valid_data(ME_L5L6_L2D4PHI3X2_CM_L5L6_L2D4PHI3X2_wr_en),
.start(VMPROJ_L5L6_L2D4PHI3X2_start),
.done(ME_L5L6_L2D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D4PHI4X1(
.number_in_vmstubin(VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1_number),
.read_add_vmstubin(VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1_read_add),
.vmstubin(VMS_L2D4PHI4X1n4_ME_L5L6_L2D4PHI4X1),
.number_in_vmprojin(VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI4X1_ME_L5L6_L2D4PHI4X1),
.matchout(ME_L5L6_L2D4PHI4X1_CM_L5L6_L2D4PHI4X1),
.valid_data(ME_L5L6_L2D4PHI4X1_CM_L5L6_L2D4PHI4X1_wr_en),
.start(VMPROJ_L5L6_L2D4PHI4X1_start),
.done(ME_L5L6_L2D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L2D4PHI4X2(
.number_in_vmstubin(VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2_number),
.read_add_vmstubin(VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2_read_add),
.vmstubin(VMS_L2D4PHI4X2n4_ME_L5L6_L2D4PHI4X2),
.number_in_vmprojin(VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2_read_add),
.vmprojin(VMPROJ_L5L6_L2D4PHI4X2_ME_L5L6_L2D4PHI4X2),
.matchout(ME_L5L6_L2D4PHI4X2_CM_L5L6_L2D4PHI4X2),
.valid_data(ME_L5L6_L2D4PHI4X2_CM_L5L6_L2D4PHI4X2_wr_en),
.start(VMPROJ_L5L6_L2D4PHI4X2_start),
.done(ME_L5L6_L2D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D3PHI1X1(
.number_in_vmstubin(VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1_number),
.read_add_vmstubin(VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1_read_add),
.vmstubin(VMS_L3D3PHI1X1n6_ME_L5L6_L3D3PHI1X1),
.number_in_vmprojin(VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI1X1_ME_L5L6_L3D3PHI1X1),
.matchout(ME_L5L6_L3D3PHI1X1_CM_L5L6_L3D3PHI1X1),
.valid_data(ME_L5L6_L3D3PHI1X1_CM_L5L6_L3D3PHI1X1_wr_en),
.start(VMPROJ_L5L6_L3D3PHI1X1_start),
.done(ME_L5L6_L3D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D3PHI1X2(
.number_in_vmstubin(VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2_number),
.read_add_vmstubin(VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2_read_add),
.vmstubin(VMS_L3D3PHI1X2n6_ME_L5L6_L3D3PHI1X2),
.number_in_vmprojin(VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI1X2_ME_L5L6_L3D3PHI1X2),
.matchout(ME_L5L6_L3D3PHI1X2_CM_L5L6_L3D3PHI1X2),
.valid_data(ME_L5L6_L3D3PHI1X2_CM_L5L6_L3D3PHI1X2_wr_en),
.start(VMPROJ_L5L6_L3D3PHI1X2_start),
.done(ME_L5L6_L3D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D3PHI2X1(
.number_in_vmstubin(VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1_number),
.read_add_vmstubin(VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1_read_add),
.vmstubin(VMS_L3D3PHI2X1n6_ME_L5L6_L3D3PHI2X1),
.number_in_vmprojin(VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI2X1_ME_L5L6_L3D3PHI2X1),
.matchout(ME_L5L6_L3D3PHI2X1_CM_L5L6_L3D3PHI2X1),
.valid_data(ME_L5L6_L3D3PHI2X1_CM_L5L6_L3D3PHI2X1_wr_en),
.start(VMPROJ_L5L6_L3D3PHI2X1_start),
.done(ME_L5L6_L3D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D3PHI2X2(
.number_in_vmstubin(VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2_number),
.read_add_vmstubin(VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2_read_add),
.vmstubin(VMS_L3D3PHI2X2n6_ME_L5L6_L3D3PHI2X2),
.number_in_vmprojin(VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI2X2_ME_L5L6_L3D3PHI2X2),
.matchout(ME_L5L6_L3D3PHI2X2_CM_L5L6_L3D3PHI2X2),
.valid_data(ME_L5L6_L3D3PHI2X2_CM_L5L6_L3D3PHI2X2_wr_en),
.start(VMPROJ_L5L6_L3D3PHI2X2_start),
.done(ME_L5L6_L3D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D3PHI3X1(
.number_in_vmstubin(VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1_number),
.read_add_vmstubin(VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1_read_add),
.vmstubin(VMS_L3D3PHI3X1n6_ME_L5L6_L3D3PHI3X1),
.number_in_vmprojin(VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI3X1_ME_L5L6_L3D3PHI3X1),
.matchout(ME_L5L6_L3D3PHI3X1_CM_L5L6_L3D3PHI3X1),
.valid_data(ME_L5L6_L3D3PHI3X1_CM_L5L6_L3D3PHI3X1_wr_en),
.start(VMPROJ_L5L6_L3D3PHI3X1_start),
.done(ME_L5L6_L3D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D3PHI3X2(
.number_in_vmstubin(VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2_number),
.read_add_vmstubin(VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2_read_add),
.vmstubin(VMS_L3D3PHI3X2n6_ME_L5L6_L3D3PHI3X2),
.number_in_vmprojin(VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2_read_add),
.vmprojin(VMPROJ_L5L6_L3D3PHI3X2_ME_L5L6_L3D3PHI3X2),
.matchout(ME_L5L6_L3D3PHI3X2_CM_L5L6_L3D3PHI3X2),
.valid_data(ME_L5L6_L3D3PHI3X2_CM_L5L6_L3D3PHI3X2_wr_en),
.start(VMPROJ_L5L6_L3D3PHI3X2_start),
.done(ME_L5L6_L3D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D4PHI1X1(
.number_in_vmstubin(VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1_number),
.read_add_vmstubin(VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1_read_add),
.vmstubin(VMS_L3D4PHI1X1n6_ME_L5L6_L3D4PHI1X1),
.number_in_vmprojin(VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI1X1_ME_L5L6_L3D4PHI1X1),
.matchout(ME_L5L6_L3D4PHI1X1_CM_L5L6_L3D4PHI1X1),
.valid_data(ME_L5L6_L3D4PHI1X1_CM_L5L6_L3D4PHI1X1_wr_en),
.start(VMPROJ_L5L6_L3D4PHI1X1_start),
.done(ME_L5L6_L3D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D4PHI1X2(
.number_in_vmstubin(VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2_number),
.read_add_vmstubin(VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2_read_add),
.vmstubin(VMS_L3D4PHI1X2n4_ME_L5L6_L3D4PHI1X2),
.number_in_vmprojin(VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI1X2_ME_L5L6_L3D4PHI1X2),
.matchout(ME_L5L6_L3D4PHI1X2_CM_L5L6_L3D4PHI1X2),
.valid_data(ME_L5L6_L3D4PHI1X2_CM_L5L6_L3D4PHI1X2_wr_en),
.start(VMPROJ_L5L6_L3D4PHI1X2_start),
.done(ME_L5L6_L3D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D4PHI2X1(
.number_in_vmstubin(VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1_number),
.read_add_vmstubin(VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1_read_add),
.vmstubin(VMS_L3D4PHI2X1n6_ME_L5L6_L3D4PHI2X1),
.number_in_vmprojin(VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI2X1_ME_L5L6_L3D4PHI2X1),
.matchout(ME_L5L6_L3D4PHI2X1_CM_L5L6_L3D4PHI2X1),
.valid_data(ME_L5L6_L3D4PHI2X1_CM_L5L6_L3D4PHI2X1_wr_en),
.start(VMPROJ_L5L6_L3D4PHI2X1_start),
.done(ME_L5L6_L3D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D4PHI2X2(
.number_in_vmstubin(VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2_number),
.read_add_vmstubin(VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2_read_add),
.vmstubin(VMS_L3D4PHI2X2n4_ME_L5L6_L3D4PHI2X2),
.number_in_vmprojin(VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI2X2_ME_L5L6_L3D4PHI2X2),
.matchout(ME_L5L6_L3D4PHI2X2_CM_L5L6_L3D4PHI2X2),
.valid_data(ME_L5L6_L3D4PHI2X2_CM_L5L6_L3D4PHI2X2_wr_en),
.start(VMPROJ_L5L6_L3D4PHI2X2_start),
.done(ME_L5L6_L3D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D4PHI3X1(
.number_in_vmstubin(VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1_number),
.read_add_vmstubin(VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1_read_add),
.vmstubin(VMS_L3D4PHI3X1n6_ME_L5L6_L3D4PHI3X1),
.number_in_vmprojin(VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI3X1_ME_L5L6_L3D4PHI3X1),
.matchout(ME_L5L6_L3D4PHI3X1_CM_L5L6_L3D4PHI3X1),
.valid_data(ME_L5L6_L3D4PHI3X1_CM_L5L6_L3D4PHI3X1_wr_en),
.start(VMPROJ_L5L6_L3D4PHI3X1_start),
.done(ME_L5L6_L3D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L3D4PHI3X2(
.number_in_vmstubin(VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2_number),
.read_add_vmstubin(VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2_read_add),
.vmstubin(VMS_L3D4PHI3X2n4_ME_L5L6_L3D4PHI3X2),
.number_in_vmprojin(VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2_read_add),
.vmprojin(VMPROJ_L5L6_L3D4PHI3X2_ME_L5L6_L3D4PHI3X2),
.matchout(ME_L5L6_L3D4PHI3X2_CM_L5L6_L3D4PHI3X2),
.valid_data(ME_L5L6_L3D4PHI3X2_CM_L5L6_L3D4PHI3X2_wr_en),
.start(VMPROJ_L5L6_L3D4PHI3X2_start),
.done(ME_L5L6_L3D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D3PHI1X1(
.number_in_vmstubin(VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1_number),
.read_add_vmstubin(VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1_read_add),
.vmstubin(VMS_L4D3PHI1X1n3_ME_L5L6_L4D3PHI1X1),
.number_in_vmprojin(VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI1X1_ME_L5L6_L4D3PHI1X1),
.matchout(ME_L5L6_L4D3PHI1X1_CM_L5L6_L4D3PHI1X1),
.valid_data(ME_L5L6_L4D3PHI1X1_CM_L5L6_L4D3PHI1X1_wr_en),
.start(VMPROJ_L5L6_L4D3PHI1X1_start),
.done(ME_L5L6_L4D3PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D3PHI1X2(
.number_in_vmstubin(VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2_number),
.read_add_vmstubin(VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2_read_add),
.vmstubin(VMS_L4D3PHI1X2n4_ME_L5L6_L4D3PHI1X2),
.number_in_vmprojin(VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI1X2_ME_L5L6_L4D3PHI1X2),
.matchout(ME_L5L6_L4D3PHI1X2_CM_L5L6_L4D3PHI1X2),
.valid_data(ME_L5L6_L4D3PHI1X2_CM_L5L6_L4D3PHI1X2_wr_en),
.start(VMPROJ_L5L6_L4D3PHI1X2_start),
.done(ME_L5L6_L4D3PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D3PHI2X1(
.number_in_vmstubin(VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1_number),
.read_add_vmstubin(VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1_read_add),
.vmstubin(VMS_L4D3PHI2X1n4_ME_L5L6_L4D3PHI2X1),
.number_in_vmprojin(VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI2X1_ME_L5L6_L4D3PHI2X1),
.matchout(ME_L5L6_L4D3PHI2X1_CM_L5L6_L4D3PHI2X1),
.valid_data(ME_L5L6_L4D3PHI2X1_CM_L5L6_L4D3PHI2X1_wr_en),
.start(VMPROJ_L5L6_L4D3PHI2X1_start),
.done(ME_L5L6_L4D3PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D3PHI2X2(
.number_in_vmstubin(VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2_number),
.read_add_vmstubin(VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2_read_add),
.vmstubin(VMS_L4D3PHI2X2n6_ME_L5L6_L4D3PHI2X2),
.number_in_vmprojin(VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI2X2_ME_L5L6_L4D3PHI2X2),
.matchout(ME_L5L6_L4D3PHI2X2_CM_L5L6_L4D3PHI2X2),
.valid_data(ME_L5L6_L4D3PHI2X2_CM_L5L6_L4D3PHI2X2_wr_en),
.start(VMPROJ_L5L6_L4D3PHI2X2_start),
.done(ME_L5L6_L4D3PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D3PHI3X1(
.number_in_vmstubin(VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1_number),
.read_add_vmstubin(VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1_read_add),
.vmstubin(VMS_L4D3PHI3X1n4_ME_L5L6_L4D3PHI3X1),
.number_in_vmprojin(VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI3X1_ME_L5L6_L4D3PHI3X1),
.matchout(ME_L5L6_L4D3PHI3X1_CM_L5L6_L4D3PHI3X1),
.valid_data(ME_L5L6_L4D3PHI3X1_CM_L5L6_L4D3PHI3X1_wr_en),
.start(VMPROJ_L5L6_L4D3PHI3X1_start),
.done(ME_L5L6_L4D3PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D3PHI3X2(
.number_in_vmstubin(VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2_number),
.read_add_vmstubin(VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2_read_add),
.vmstubin(VMS_L4D3PHI3X2n6_ME_L5L6_L4D3PHI3X2),
.number_in_vmprojin(VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI3X2_ME_L5L6_L4D3PHI3X2),
.matchout(ME_L5L6_L4D3PHI3X2_CM_L5L6_L4D3PHI3X2),
.valid_data(ME_L5L6_L4D3PHI3X2_CM_L5L6_L4D3PHI3X2_wr_en),
.start(VMPROJ_L5L6_L4D3PHI3X2_start),
.done(ME_L5L6_L4D3PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D3PHI4X1(
.number_in_vmstubin(VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1_number),
.read_add_vmstubin(VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1_read_add),
.vmstubin(VMS_L4D3PHI4X1n3_ME_L5L6_L4D3PHI4X1),
.number_in_vmprojin(VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI4X1_ME_L5L6_L4D3PHI4X1),
.matchout(ME_L5L6_L4D3PHI4X1_CM_L5L6_L4D3PHI4X1),
.valid_data(ME_L5L6_L4D3PHI4X1_CM_L5L6_L4D3PHI4X1_wr_en),
.start(VMPROJ_L5L6_L4D3PHI4X1_start),
.done(ME_L5L6_L4D3PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D3PHI4X2(
.number_in_vmstubin(VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2_number),
.read_add_vmstubin(VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2_read_add),
.vmstubin(VMS_L4D3PHI4X2n4_ME_L5L6_L4D3PHI4X2),
.number_in_vmprojin(VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2_read_add),
.vmprojin(VMPROJ_L5L6_L4D3PHI4X2_ME_L5L6_L4D3PHI4X2),
.matchout(ME_L5L6_L4D3PHI4X2_CM_L5L6_L4D3PHI4X2),
.valid_data(ME_L5L6_L4D3PHI4X2_CM_L5L6_L4D3PHI4X2_wr_en),
.start(VMPROJ_L5L6_L4D3PHI4X2_start),
.done(ME_L5L6_L4D3PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D4PHI1X1(
.number_in_vmstubin(VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1_number),
.read_add_vmstubin(VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1_read_add),
.vmstubin(VMS_L4D4PHI1X1n4_ME_L5L6_L4D4PHI1X1),
.number_in_vmprojin(VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI1X1_ME_L5L6_L4D4PHI1X1),
.matchout(ME_L5L6_L4D4PHI1X1_CM_L5L6_L4D4PHI1X1),
.valid_data(ME_L5L6_L4D4PHI1X1_CM_L5L6_L4D4PHI1X1_wr_en),
.start(VMPROJ_L5L6_L4D4PHI1X1_start),
.done(ME_L5L6_L4D4PHI1X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D4PHI1X2(
.number_in_vmstubin(VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2_number),
.read_add_vmstubin(VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2_read_add),
.vmstubin(VMS_L4D4PHI1X2n4_ME_L5L6_L4D4PHI1X2),
.number_in_vmprojin(VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI1X2_ME_L5L6_L4D4PHI1X2),
.matchout(ME_L5L6_L4D4PHI1X2_CM_L5L6_L4D4PHI1X2),
.valid_data(ME_L5L6_L4D4PHI1X2_CM_L5L6_L4D4PHI1X2_wr_en),
.start(VMPROJ_L5L6_L4D4PHI1X2_start),
.done(ME_L5L6_L4D4PHI1X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D4PHI2X1(
.number_in_vmstubin(VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1_number),
.read_add_vmstubin(VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1_read_add),
.vmstubin(VMS_L4D4PHI2X1n6_ME_L5L6_L4D4PHI2X1),
.number_in_vmprojin(VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI2X1_ME_L5L6_L4D4PHI2X1),
.matchout(ME_L5L6_L4D4PHI2X1_CM_L5L6_L4D4PHI2X1),
.valid_data(ME_L5L6_L4D4PHI2X1_CM_L5L6_L4D4PHI2X1_wr_en),
.start(VMPROJ_L5L6_L4D4PHI2X1_start),
.done(ME_L5L6_L4D4PHI2X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D4PHI2X2(
.number_in_vmstubin(VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2_number),
.read_add_vmstubin(VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2_read_add),
.vmstubin(VMS_L4D4PHI2X2n6_ME_L5L6_L4D4PHI2X2),
.number_in_vmprojin(VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI2X2_ME_L5L6_L4D4PHI2X2),
.matchout(ME_L5L6_L4D4PHI2X2_CM_L5L6_L4D4PHI2X2),
.valid_data(ME_L5L6_L4D4PHI2X2_CM_L5L6_L4D4PHI2X2_wr_en),
.start(VMPROJ_L5L6_L4D4PHI2X2_start),
.done(ME_L5L6_L4D4PHI2X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D4PHI3X1(
.number_in_vmstubin(VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1_number),
.read_add_vmstubin(VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1_read_add),
.vmstubin(VMS_L4D4PHI3X1n6_ME_L5L6_L4D4PHI3X1),
.number_in_vmprojin(VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI3X1_ME_L5L6_L4D4PHI3X1),
.matchout(ME_L5L6_L4D4PHI3X1_CM_L5L6_L4D4PHI3X1),
.valid_data(ME_L5L6_L4D4PHI3X1_CM_L5L6_L4D4PHI3X1_wr_en),
.start(VMPROJ_L5L6_L4D4PHI3X1_start),
.done(ME_L5L6_L4D4PHI3X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D4PHI3X2(
.number_in_vmstubin(VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2_number),
.read_add_vmstubin(VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2_read_add),
.vmstubin(VMS_L4D4PHI3X2n6_ME_L5L6_L4D4PHI3X2),
.number_in_vmprojin(VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI3X2_ME_L5L6_L4D4PHI3X2),
.matchout(ME_L5L6_L4D4PHI3X2_CM_L5L6_L4D4PHI3X2),
.valid_data(ME_L5L6_L4D4PHI3X2_CM_L5L6_L4D4PHI3X2_wr_en),
.start(VMPROJ_L5L6_L4D4PHI3X2_start),
.done(ME_L5L6_L4D4PHI3X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D4PHI4X1(
.number_in_vmstubin(VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1_number),
.read_add_vmstubin(VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1_read_add),
.vmstubin(VMS_L4D4PHI4X1n4_ME_L5L6_L4D4PHI4X1),
.number_in_vmprojin(VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI4X1_ME_L5L6_L4D4PHI4X1),
.matchout(ME_L5L6_L4D4PHI4X1_CM_L5L6_L4D4PHI4X1),
.valid_data(ME_L5L6_L4D4PHI4X1_CM_L5L6_L4D4PHI4X1_wr_en),
.start(VMPROJ_L5L6_L4D4PHI4X1_start),
.done(ME_L5L6_L4D4PHI4X1_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchEngine  ME_L5L6_L4D4PHI4X2(
.number_in_vmstubin(VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2_number),
.read_add_vmstubin(VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2_read_add),
.vmstubin(VMS_L4D4PHI4X2n4_ME_L5L6_L4D4PHI4X2),
.number_in_vmprojin(VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2_number),
.read_add_vmprojin(VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2_read_add),
.vmprojin(VMPROJ_L5L6_L4D4PHI4X2_ME_L5L6_L4D4PHI4X2),
.matchout(ME_L5L6_L4D4PHI4X2_CM_L5L6_L4D4PHI4X2),
.valid_data(ME_L5L6_L4D4PHI4X2_CM_L5L6_L4D4PHI4X2_wr_en),
.start(VMPROJ_L5L6_L4D4PHI4X2_start),
.done(ME_L5L6_L4D4PHI4X2_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b1,`PHI_L1,`Z_L1,`R_L1,`PHID_L1,`ZD_L1,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L3L4_L1,`MC_z_L3L4_L1,`MC_zfactor_INNER) MC_L3L4_L1D3(
.number_in_match1in(CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3_number),
.read_add_match1in(CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3_read_add),
.match1in(CM_L3L4_L1D3PHI1X1_MC_L3L4_L1D3),
.number_in_match2in(CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3_number),
.read_add_match2in(CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3_read_add),
.match2in(CM_L3L4_L1D3PHI1X2_MC_L3L4_L1D3),
.number_in_match3in(CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3_number),
.read_add_match3in(CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3_read_add),
.match3in(CM_L3L4_L1D3PHI2X1_MC_L3L4_L1D3),
.number_in_match4in(CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3_number),
.read_add_match4in(CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3_read_add),
.match4in(CM_L3L4_L1D3PHI2X2_MC_L3L4_L1D3),
.number_in_match5in(CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3_number),
.read_add_match5in(CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3_read_add),
.match5in(CM_L3L4_L1D3PHI3X1_MC_L3L4_L1D3),
.number_in_match6in(CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3_number),
.read_add_match6in(CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3_read_add),
.match6in(CM_L3L4_L1D3PHI3X2_MC_L3L4_L1D3),
.read_add_allprojin(AP_L3L4_L1D3_MC_L3L4_L1D3_read_add),
.allprojin(AP_L3L4_L1D3_MC_L3L4_L1D3),
.read_add_allstubin(AS_L1D3n3_MC_L3L4_L1D3_read_add),
.allstubin(AS_L1D3n3_MC_L3L4_L1D3),
.matchoutminus(MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus),
.matchoutplus(MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus),
.matchout1(MC_L3L4_L1D3_FM_L3L4_L1D3),
.valid_matchminus(MC_L3L4_L1D3_FM_L3L4_L1D3_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L1D3_FM_L3L4_L1D3_ToPlus_wr_en),
.valid_match(MC_L3L4_L1D3_FM_L3L4_L1D3_wr_en),
.start(CM_L3L4_L1D3PHI1X1_start),
.done(MC_L3L4_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b1,`PHI_L1,`Z_L1,`R_L1,`PHID_L1,`ZD_L1,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L3L4_L1,`MC_z_L3L4_L1,`MC_zfactor_INNER) MC_L3L4_L1D4(
.number_in_match1in(CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4_number),
.read_add_match1in(CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4_read_add),
.match1in(CM_L3L4_L1D4PHI1X1_MC_L3L4_L1D4),
.number_in_match2in(CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4_number),
.read_add_match2in(CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4_read_add),
.match2in(CM_L3L4_L1D4PHI1X2_MC_L3L4_L1D4),
.number_in_match3in(CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4_number),
.read_add_match3in(CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4_read_add),
.match3in(CM_L3L4_L1D4PHI2X1_MC_L3L4_L1D4),
.number_in_match4in(CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4_number),
.read_add_match4in(CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4_read_add),
.match4in(CM_L3L4_L1D4PHI2X2_MC_L3L4_L1D4),
.number_in_match5in(CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4_number),
.read_add_match5in(CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4_read_add),
.match5in(CM_L3L4_L1D4PHI3X1_MC_L3L4_L1D4),
.number_in_match6in(CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4_number),
.read_add_match6in(CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4_read_add),
.match6in(CM_L3L4_L1D4PHI3X2_MC_L3L4_L1D4),
.read_add_allprojin(AP_L3L4_L1D4_MC_L3L4_L1D4_read_add),
.allprojin(AP_L3L4_L1D4_MC_L3L4_L1D4),
.read_add_allstubin(AS_L1D4n2_MC_L3L4_L1D4_read_add),
.allstubin(AS_L1D4n2_MC_L3L4_L1D4),
.matchoutminus(MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus),
.matchoutplus(MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus),
.matchout1(MC_L3L4_L1D4_FM_L3L4_L1D4),
.valid_matchminus(MC_L3L4_L1D4_FM_L3L4_L1D4_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L1D4_FM_L3L4_L1D4_ToPlus_wr_en),
.valid_match(MC_L3L4_L1D4_FM_L3L4_L1D4_wr_en),
.start(CM_L3L4_L1D4PHI1X1_start),
.done(MC_L3L4_L1D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b1,`PHI_L2,`Z_L2,`R_L2,`PHID_L2,`ZD_L2,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L3L4_L2,`MC_z_L3L4_L2,`MC_zfactor_INNER) MC_L3L4_L2D3(
.number_in_match1in(CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3_number),
.read_add_match1in(CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3_read_add),
.match1in(CM_L3L4_L2D3PHI1X1_MC_L3L4_L2D3),
.number_in_match2in(CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3_number),
.read_add_match2in(CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3_read_add),
.match2in(CM_L3L4_L2D3PHI1X2_MC_L3L4_L2D3),
.number_in_match3in(CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3_number),
.read_add_match3in(CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3_read_add),
.match3in(CM_L3L4_L2D3PHI2X1_MC_L3L4_L2D3),
.number_in_match4in(CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3_number),
.read_add_match4in(CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3_read_add),
.match4in(CM_L3L4_L2D3PHI2X2_MC_L3L4_L2D3),
.number_in_match5in(CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3_number),
.read_add_match5in(CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3_read_add),
.match5in(CM_L3L4_L2D3PHI3X1_MC_L3L4_L2D3),
.number_in_match6in(CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3_number),
.read_add_match6in(CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3_read_add),
.match6in(CM_L3L4_L2D3PHI3X2_MC_L3L4_L2D3),
.number_in_match7in(CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3_number),
.read_add_match7in(CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3_read_add),
.match7in(CM_L3L4_L2D3PHI4X1_MC_L3L4_L2D3),
.number_in_match8in(CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3_number),
.read_add_match8in(CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3_read_add),
.match8in(CM_L3L4_L2D3PHI4X2_MC_L3L4_L2D3),
.read_add_allprojin(AP_L3L4_L2D3_MC_L3L4_L2D3_read_add),
.allprojin(AP_L3L4_L2D3_MC_L3L4_L2D3),
.read_add_allstubin(AS_L2D3n2_MC_L3L4_L2D3_read_add),
.allstubin(AS_L2D3n2_MC_L3L4_L2D3),
.matchoutminus(MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus),
.matchoutplus(MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus),
.matchout1(MC_L3L4_L2D3_FM_L3L4_L2D3),
.valid_matchminus(MC_L3L4_L2D3_FM_L3L4_L2D3_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L2D3_FM_L3L4_L2D3_ToPlus_wr_en),
.valid_match(MC_L3L4_L2D3_FM_L3L4_L2D3_wr_en),
.start(CM_L3L4_L2D3PHI1X1_start),
.done(MC_L3L4_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b1,`PHI_L2,`Z_L2,`R_L2,`PHID_L2,`ZD_L2,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L3L4_L2,`MC_z_L3L4_L2,`MC_zfactor_INNER) MC_L3L4_L2D4(
.number_in_match1in(CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4_number),
.read_add_match1in(CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4_read_add),
.match1in(CM_L3L4_L2D4PHI1X1_MC_L3L4_L2D4),
.number_in_match2in(CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4_number),
.read_add_match2in(CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4_read_add),
.match2in(CM_L3L4_L2D4PHI1X2_MC_L3L4_L2D4),
.number_in_match3in(CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4_number),
.read_add_match3in(CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4_read_add),
.match3in(CM_L3L4_L2D4PHI2X1_MC_L3L4_L2D4),
.number_in_match4in(CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4_number),
.read_add_match4in(CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4_read_add),
.match4in(CM_L3L4_L2D4PHI2X2_MC_L3L4_L2D4),
.number_in_match5in(CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4_number),
.read_add_match5in(CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4_read_add),
.match5in(CM_L3L4_L2D4PHI3X1_MC_L3L4_L2D4),
.number_in_match6in(CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4_number),
.read_add_match6in(CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4_read_add),
.match6in(CM_L3L4_L2D4PHI3X2_MC_L3L4_L2D4),
.number_in_match7in(CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4_number),
.read_add_match7in(CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4_read_add),
.match7in(CM_L3L4_L2D4PHI4X1_MC_L3L4_L2D4),
.number_in_match8in(CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4_number),
.read_add_match8in(CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4_read_add),
.match8in(CM_L3L4_L2D4PHI4X2_MC_L3L4_L2D4),
.read_add_allprojin(AP_L3L4_L2D4_MC_L3L4_L2D4_read_add),
.allprojin(AP_L3L4_L2D4_MC_L3L4_L2D4),
.read_add_allstubin(AS_L2D4n3_MC_L3L4_L2D4_read_add),
.allstubin(AS_L2D4n3_MC_L3L4_L2D4),
.matchoutminus(MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus),
.matchoutplus(MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus),
.matchout1(MC_L3L4_L2D4_FM_L3L4_L2D4),
.valid_matchminus(MC_L3L4_L2D4_FM_L3L4_L2D4_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L2D4_FM_L3L4_L2D4_ToPlus_wr_en),
.valid_match(MC_L3L4_L2D4_FM_L3L4_L2D4_wr_en),
.start(CM_L3L4_L2D4PHI1X1_start),
.done(MC_L3L4_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b0,`PHI_L5,`Z_L5,`R_L5,`PHID_L5,`ZD_L5,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L3L4_L5,`MC_z_L3L4_L5,`MC_zfactor_OUTER) MC_L3L4_L5D3(
.number_in_match1in(CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3_number),
.read_add_match1in(CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3_read_add),
.match1in(CM_L3L4_L5D3PHI1X1_MC_L3L4_L5D3),
.number_in_match2in(CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3_number),
.read_add_match2in(CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3_read_add),
.match2in(CM_L3L4_L5D3PHI1X2_MC_L3L4_L5D3),
.number_in_match3in(CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3_number),
.read_add_match3in(CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3_read_add),
.match3in(CM_L3L4_L5D3PHI2X1_MC_L3L4_L5D3),
.number_in_match4in(CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3_number),
.read_add_match4in(CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3_read_add),
.match4in(CM_L3L4_L5D3PHI2X2_MC_L3L4_L5D3),
.number_in_match5in(CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3_number),
.read_add_match5in(CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3_read_add),
.match5in(CM_L3L4_L5D3PHI3X1_MC_L3L4_L5D3),
.number_in_match6in(CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3_number),
.read_add_match6in(CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3_read_add),
.match6in(CM_L3L4_L5D3PHI3X2_MC_L3L4_L5D3),
.read_add_allprojin(AP_L3L4_L5D3_MC_L3L4_L5D3_read_add),
.allprojin(AP_L3L4_L5D3_MC_L3L4_L5D3),
.read_add_allstubin(AS_L5D3n3_MC_L3L4_L5D3_read_add),
.allstubin(AS_L5D3n3_MC_L3L4_L5D3),
.matchoutminus(MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus),
.matchoutplus(MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus),
.matchout1(MC_L3L4_L5D3_FM_L3L4_L5D3),
.valid_matchminus(MC_L3L4_L5D3_FM_L3L4_L5D3_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L5D3_FM_L3L4_L5D3_ToPlus_wr_en),
.valid_match(MC_L3L4_L5D3_FM_L3L4_L5D3_wr_en),
.start(CM_L3L4_L5D3PHI1X1_start),
.done(MC_L3L4_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b0,`PHI_L5,`Z_L5,`R_L5,`PHID_L5,`ZD_L5,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L3L4_L5,`MC_z_L3L4_L5,`MC_zfactor_OUTER) MC_L3L4_L5D4(
.number_in_match1in(CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4_number),
.read_add_match1in(CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4_read_add),
.match1in(CM_L3L4_L5D4PHI1X1_MC_L3L4_L5D4),
.number_in_match2in(CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4_number),
.read_add_match2in(CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4_read_add),
.match2in(CM_L3L4_L5D4PHI1X2_MC_L3L4_L5D4),
.number_in_match3in(CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4_number),
.read_add_match3in(CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4_read_add),
.match3in(CM_L3L4_L5D4PHI2X1_MC_L3L4_L5D4),
.number_in_match4in(CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4_number),
.read_add_match4in(CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4_read_add),
.match4in(CM_L3L4_L5D4PHI2X2_MC_L3L4_L5D4),
.number_in_match5in(CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4_number),
.read_add_match5in(CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4_read_add),
.match5in(CM_L3L4_L5D4PHI3X1_MC_L3L4_L5D4),
.number_in_match6in(CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4_number),
.read_add_match6in(CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4_read_add),
.match6in(CM_L3L4_L5D4PHI3X2_MC_L3L4_L5D4),
.read_add_allprojin(AP_L3L4_L5D4_MC_L3L4_L5D4_read_add),
.allprojin(AP_L3L4_L5D4_MC_L3L4_L5D4),
.read_add_allstubin(AS_L5D4n2_MC_L3L4_L5D4_read_add),
.allstubin(AS_L5D4n2_MC_L3L4_L5D4),
.matchoutminus(MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus),
.matchoutplus(MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus),
.matchout1(MC_L3L4_L5D4_FM_L3L4_L5D4),
.valid_matchminus(MC_L3L4_L5D4_FM_L3L4_L5D4_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L5D4_FM_L3L4_L5D4_ToPlus_wr_en),
.valid_match(MC_L3L4_L5D4_FM_L3L4_L5D4_wr_en),
.start(CM_L3L4_L5D4PHI1X1_start),
.done(MC_L3L4_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b0,`PHI_L6,`Z_L6,`R_L6,`PHID_L6,`ZD_L6,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L3L4_L6,`MC_z_L3L4_L6,`MC_zfactor_OUTER) MC_L3L4_L6D3(
.number_in_match1in(CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3_number),
.read_add_match1in(CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3_read_add),
.match1in(CM_L3L4_L6D3PHI1X1_MC_L3L4_L6D3),
.number_in_match2in(CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3_number),
.read_add_match2in(CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3_read_add),
.match2in(CM_L3L4_L6D3PHI1X2_MC_L3L4_L6D3),
.number_in_match3in(CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3_number),
.read_add_match3in(CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3_read_add),
.match3in(CM_L3L4_L6D3PHI2X1_MC_L3L4_L6D3),
.number_in_match4in(CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3_number),
.read_add_match4in(CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3_read_add),
.match4in(CM_L3L4_L6D3PHI2X2_MC_L3L4_L6D3),
.number_in_match5in(CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3_number),
.read_add_match5in(CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3_read_add),
.match5in(CM_L3L4_L6D3PHI3X1_MC_L3L4_L6D3),
.number_in_match6in(CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3_number),
.read_add_match6in(CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3_read_add),
.match6in(CM_L3L4_L6D3PHI3X2_MC_L3L4_L6D3),
.number_in_match7in(CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3_number),
.read_add_match7in(CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3_read_add),
.match7in(CM_L3L4_L6D3PHI4X1_MC_L3L4_L6D3),
.number_in_match8in(CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3_number),
.read_add_match8in(CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3_read_add),
.match8in(CM_L3L4_L6D3PHI4X2_MC_L3L4_L6D3),
.read_add_allprojin(AP_L3L4_L6D3_MC_L3L4_L6D3_read_add),
.allprojin(AP_L3L4_L6D3_MC_L3L4_L6D3),
.read_add_allstubin(AS_L6D3n2_MC_L3L4_L6D3_read_add),
.allstubin(AS_L6D3n2_MC_L3L4_L6D3),
.matchoutminus(MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus),
.matchoutplus(MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus),
.matchout1(MC_L3L4_L6D3_FM_L3L4_L6D3),
.valid_matchminus(MC_L3L4_L6D3_FM_L3L4_L6D3_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L6D3_FM_L3L4_L6D3_ToPlus_wr_en),
.valid_match(MC_L3L4_L6D3_FM_L3L4_L6D3_wr_en),
.start(CM_L3L4_L6D3PHI1X1_start),
.done(MC_L3L4_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b0,`PHI_L6,`Z_L6,`R_L6,`PHID_L6,`ZD_L6,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L3L4_L6,`MC_z_L3L4_L6,`MC_zfactor_OUTER) MC_L3L4_L6D4(
.number_in_match1in(CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4_number),
.read_add_match1in(CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4_read_add),
.match1in(CM_L3L4_L6D4PHI1X1_MC_L3L4_L6D4),
.number_in_match2in(CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4_number),
.read_add_match2in(CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4_read_add),
.match2in(CM_L3L4_L6D4PHI1X2_MC_L3L4_L6D4),
.number_in_match3in(CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4_number),
.read_add_match3in(CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4_read_add),
.match3in(CM_L3L4_L6D4PHI2X1_MC_L3L4_L6D4),
.number_in_match4in(CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4_number),
.read_add_match4in(CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4_read_add),
.match4in(CM_L3L4_L6D4PHI2X2_MC_L3L4_L6D4),
.number_in_match5in(CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4_number),
.read_add_match5in(CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4_read_add),
.match5in(CM_L3L4_L6D4PHI3X1_MC_L3L4_L6D4),
.number_in_match6in(CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4_number),
.read_add_match6in(CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4_read_add),
.match6in(CM_L3L4_L6D4PHI3X2_MC_L3L4_L6D4),
.number_in_match7in(CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4_number),
.read_add_match7in(CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4_read_add),
.match7in(CM_L3L4_L6D4PHI4X1_MC_L3L4_L6D4),
.number_in_match8in(CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4_number),
.read_add_match8in(CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4_read_add),
.match8in(CM_L3L4_L6D4PHI4X2_MC_L3L4_L6D4),
.read_add_allprojin(AP_L3L4_L6D4_MC_L3L4_L6D4_read_add),
.allprojin(AP_L3L4_L6D4_MC_L3L4_L6D4),
.read_add_allstubin(AS_L6D4n3_MC_L3L4_L6D4_read_add),
.allstubin(AS_L6D4n3_MC_L3L4_L6D4),
.matchoutminus(MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus),
.matchoutplus(MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus),
.matchout1(MC_L3L4_L6D4_FM_L3L4_L6D4),
.valid_matchminus(MC_L3L4_L6D4_FM_L3L4_L6D4_ToMinus_wr_en),
.valid_matchplus(MC_L3L4_L6D4_FM_L3L4_L6D4_ToPlus_wr_en),
.valid_match(MC_L3L4_L6D4_FM_L3L4_L6D4_wr_en),
.start(CM_L3L4_L6D4PHI1X1_start),
.done(MC_L3L4_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b1,`PHI_L1,`Z_L1,`R_L1,`PHID_L1,`ZD_L1,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L1,`MC_z_L5L6_L1,`MC_zfactor_INNER) MC_L5L6_L1D3(
.number_in_match1in(CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3_number),
.read_add_match1in(CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3_read_add),
.match1in(CM_L5L6_L1D3PHI1X1_MC_L5L6_L1D3),
.number_in_match2in(CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3_number),
.read_add_match2in(CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3_read_add),
.match2in(CM_L5L6_L1D3PHI1X2_MC_L5L6_L1D3),
.number_in_match3in(CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3_number),
.read_add_match3in(CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3_read_add),
.match3in(CM_L5L6_L1D3PHI2X1_MC_L5L6_L1D3),
.number_in_match4in(CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3_number),
.read_add_match4in(CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3_read_add),
.match4in(CM_L5L6_L1D3PHI2X2_MC_L5L6_L1D3),
.number_in_match5in(CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3_number),
.read_add_match5in(CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3_read_add),
.match5in(CM_L5L6_L1D3PHI3X1_MC_L5L6_L1D3),
.number_in_match6in(CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3_number),
.read_add_match6in(CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3_read_add),
.match6in(CM_L5L6_L1D3PHI3X2_MC_L5L6_L1D3),
.read_add_allprojin(AP_L5L6_L1D3_MC_L5L6_L1D3_read_add),
.allprojin(AP_L5L6_L1D3_MC_L5L6_L1D3),
.read_add_allstubin(AS_L1D3n4_MC_L5L6_L1D3_read_add),
.allstubin(AS_L1D3n4_MC_L5L6_L1D3),
.matchoutminus(MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus),
.matchoutplus(MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus),
.matchout1(MC_L5L6_L1D3_FM_L5L6_L1D3),
.valid_matchminus(MC_L5L6_L1D3_FM_L5L6_L1D3_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L1D3_FM_L5L6_L1D3_ToPlus_wr_en),
.valid_match(MC_L5L6_L1D3_FM_L5L6_L1D3_wr_en),
.start(CM_L5L6_L1D3PHI1X1_start),
.done(MC_L5L6_L1D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b1,`PHI_L1,`Z_L1,`R_L1,`PHID_L1,`ZD_L1,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L1,`MC_z_L5L6_L1,`MC_zfactor_INNER) MC_L5L6_L1D4(
.number_in_match1in(CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4_number),
.read_add_match1in(CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4_read_add),
.match1in(CM_L5L6_L1D4PHI1X1_MC_L5L6_L1D4),
.number_in_match2in(CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4_number),
.read_add_match2in(CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4_read_add),
.match2in(CM_L5L6_L1D4PHI1X2_MC_L5L6_L1D4),
.number_in_match3in(CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4_number),
.read_add_match3in(CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4_read_add),
.match3in(CM_L5L6_L1D4PHI2X1_MC_L5L6_L1D4),
.number_in_match4in(CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4_number),
.read_add_match4in(CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4_read_add),
.match4in(CM_L5L6_L1D4PHI2X2_MC_L5L6_L1D4),
.number_in_match5in(CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4_number),
.read_add_match5in(CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4_read_add),
.match5in(CM_L5L6_L1D4PHI3X1_MC_L5L6_L1D4),
.number_in_match6in(CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4_number),
.read_add_match6in(CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4_read_add),
.match6in(CM_L5L6_L1D4PHI3X2_MC_L5L6_L1D4),
.read_add_allprojin(AP_L5L6_L1D4_MC_L5L6_L1D4_read_add),
.allprojin(AP_L5L6_L1D4_MC_L5L6_L1D4),
.read_add_allstubin(AS_L1D4n3_MC_L5L6_L1D4_read_add),
.allstubin(AS_L1D4n3_MC_L5L6_L1D4),
.matchoutminus(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus),
.matchoutplus(MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus),
.matchout1(MC_L5L6_L1D4_FM_L5L6_L1D4),
.valid_matchminus(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L1D4_FM_L5L6_L1D4_ToPlus_wr_en),
.valid_match(MC_L5L6_L1D4_FM_L5L6_L1D4_wr_en),
.valid_match2(MC_L5L6_L1D4_FM_L5L6_L1D4_ToMinus_wr_en_wr_en),
.start(CM_L5L6_L1D4PHI1X1_start),
.done(MC_L5L6_L1D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b1,`PHI_L2,`Z_L2,`R_L2,`PHID_L2,`ZD_L2,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L2,`MC_z_L5L6_L2,`MC_zfactor_INNER) MC_L5L6_L2D3(
.number_in_match1in(CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3_number),
.read_add_match1in(CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3_read_add),
.match1in(CM_L5L6_L2D3PHI1X1_MC_L5L6_L2D3),
.number_in_match2in(CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3_number),
.read_add_match2in(CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3_read_add),
.match2in(CM_L5L6_L2D3PHI1X2_MC_L5L6_L2D3),
.number_in_match3in(CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3_number),
.read_add_match3in(CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3_read_add),
.match3in(CM_L5L6_L2D3PHI2X1_MC_L5L6_L2D3),
.number_in_match4in(CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3_number),
.read_add_match4in(CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3_read_add),
.match4in(CM_L5L6_L2D3PHI2X2_MC_L5L6_L2D3),
.number_in_match5in(CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3_number),
.read_add_match5in(CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3_read_add),
.match5in(CM_L5L6_L2D3PHI3X1_MC_L5L6_L2D3),
.number_in_match6in(CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3_number),
.read_add_match6in(CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3_read_add),
.match6in(CM_L5L6_L2D3PHI3X2_MC_L5L6_L2D3),
.number_in_match7in(CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3_number),
.read_add_match7in(CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3_read_add),
.match7in(CM_L5L6_L2D3PHI4X1_MC_L5L6_L2D3),
.number_in_match8in(CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3_number),
.read_add_match8in(CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3_read_add),
.match8in(CM_L5L6_L2D3PHI4X2_MC_L5L6_L2D3),
.read_add_allprojin(AP_L5L6_L2D3_MC_L5L6_L2D3_read_add),
.allprojin(AP_L5L6_L2D3_MC_L5L6_L2D3),
.read_add_allstubin(AS_L2D3n3_MC_L5L6_L2D3_read_add),
.allstubin(AS_L2D3n3_MC_L5L6_L2D3),
.matchoutminus(MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus),
.matchoutplus(MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus),
.matchout1(MC_L5L6_L2D3_FM_L5L6_L2D3),
.valid_matchminus(MC_L5L6_L2D3_FM_L5L6_L2D3_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L2D3_FM_L5L6_L2D3_ToPlus_wr_en),
.valid_match(MC_L5L6_L2D3_FM_L5L6_L2D3_wr_en),
.start(CM_L5L6_L2D3PHI1X1_start),
.done(MC_L5L6_L2D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b1,`PHI_L2,`Z_L2,`R_L2,`PHID_L2,`ZD_L2,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L2,`MC_z_L5L6_L2,`MC_zfactor_INNER) MC_L5L6_L2D4(
.number_in_match1in(CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4_number),
.read_add_match1in(CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4_read_add),
.match1in(CM_L5L6_L2D4PHI1X1_MC_L5L6_L2D4),
.number_in_match2in(CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4_number),
.read_add_match2in(CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4_read_add),
.match2in(CM_L5L6_L2D4PHI1X2_MC_L5L6_L2D4),
.number_in_match3in(CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4_number),
.read_add_match3in(CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4_read_add),
.match3in(CM_L5L6_L2D4PHI2X1_MC_L5L6_L2D4),
.number_in_match4in(CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4_number),
.read_add_match4in(CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4_read_add),
.match4in(CM_L5L6_L2D4PHI2X2_MC_L5L6_L2D4),
.number_in_match5in(CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4_number),
.read_add_match5in(CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4_read_add),
.match5in(CM_L5L6_L2D4PHI3X1_MC_L5L6_L2D4),
.number_in_match6in(CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4_number),
.read_add_match6in(CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4_read_add),
.match6in(CM_L5L6_L2D4PHI3X2_MC_L5L6_L2D4),
.number_in_match7in(CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4_number),
.read_add_match7in(CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4_read_add),
.match7in(CM_L5L6_L2D4PHI4X1_MC_L5L6_L2D4),
.number_in_match8in(CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4_number),
.read_add_match8in(CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4_read_add),
.match8in(CM_L5L6_L2D4PHI4X2_MC_L5L6_L2D4),
.read_add_allprojin(AP_L5L6_L2D4_MC_L5L6_L2D4_read_add),
.allprojin(AP_L5L6_L2D4_MC_L5L6_L2D4),
.read_add_allstubin(AS_L2D4n4_MC_L5L6_L2D4_read_add),
.allstubin(AS_L2D4n4_MC_L5L6_L2D4),
.matchoutminus(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus),
.matchoutplus(MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus),
.matchout1(MC_L5L6_L2D4_FM_L5L6_L2D4),
.valid_matchminus(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L2D4_FM_L5L6_L2D4_ToPlus_wr_en),
.valid_match(MC_L5L6_L2D4_FM_L5L6_L2D4_wr_en),
.valid_match2(MC_L5L6_L2D4_FM_L5L6_L2D4_ToMinus_wr_en_wr_en),
.start(CM_L5L6_L2D4PHI1X1_start),
.done(MC_L5L6_L2D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b1,`PHI_L3,`Z_L3,`R_L3,`PHID_L3,`ZD_L3,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L3,`MC_z_L5L6_L3,`MC_zfactor_INNER) MC_L5L6_L3D3(
.number_in_match1in(CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3_number),
.read_add_match1in(CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3_read_add),
.match1in(CM_L5L6_L3D3PHI1X1_MC_L5L6_L3D3),
.number_in_match2in(CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3_number),
.read_add_match2in(CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3_read_add),
.match2in(CM_L5L6_L3D3PHI1X2_MC_L5L6_L3D3),
.number_in_match3in(CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3_number),
.read_add_match3in(CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3_read_add),
.match3in(CM_L5L6_L3D3PHI2X1_MC_L5L6_L3D3),
.number_in_match4in(CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3_number),
.read_add_match4in(CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3_read_add),
.match4in(CM_L5L6_L3D3PHI2X2_MC_L5L6_L3D3),
.number_in_match5in(CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3_number),
.read_add_match5in(CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3_read_add),
.match5in(CM_L5L6_L3D3PHI3X1_MC_L5L6_L3D3),
.number_in_match6in(CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3_number),
.read_add_match6in(CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3_read_add),
.match6in(CM_L5L6_L3D3PHI3X2_MC_L5L6_L3D3),
.read_add_allprojin(AP_L5L6_L3D3_MC_L5L6_L3D3_read_add),
.allprojin(AP_L5L6_L3D3_MC_L5L6_L3D3),
.read_add_allstubin(AS_L3D3n3_MC_L5L6_L3D3_read_add),
.allstubin(AS_L3D3n3_MC_L5L6_L3D3),
.matchoutminus(MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus),
.matchoutplus(MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus),
.matchout1(MC_L5L6_L3D3_FM_L5L6_L3D3),
.valid_matchminus(MC_L5L6_L3D3_FM_L5L6_L3D3_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L3D3_FM_L5L6_L3D3_ToPlus_wr_en),
.valid_match(MC_L5L6_L3D3_FM_L5L6_L3D3_wr_en),
.start(CM_L5L6_L3D3PHI1X1_start),
.done(MC_L5L6_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b1,`PHI_L3,`Z_L3,`R_L3,`PHID_L3,`ZD_L3,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L5L6_L3,`MC_z_L5L6_L3,`MC_zfactor_INNER) MC_L5L6_L3D4(
.number_in_match1in(CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4_number),
.read_add_match1in(CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4_read_add),
.match1in(CM_L5L6_L3D4PHI1X1_MC_L5L6_L3D4),
.number_in_match2in(CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4_number),
.read_add_match2in(CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4_read_add),
.match2in(CM_L5L6_L3D4PHI1X2_MC_L5L6_L3D4),
.number_in_match3in(CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4_number),
.read_add_match3in(CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4_read_add),
.match3in(CM_L5L6_L3D4PHI2X1_MC_L5L6_L3D4),
.number_in_match4in(CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4_number),
.read_add_match4in(CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4_read_add),
.match4in(CM_L5L6_L3D4PHI2X2_MC_L5L6_L3D4),
.number_in_match5in(CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4_number),
.read_add_match5in(CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4_read_add),
.match5in(CM_L5L6_L3D4PHI3X1_MC_L5L6_L3D4),
.number_in_match6in(CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4_number),
.read_add_match6in(CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4_read_add),
.match6in(CM_L5L6_L3D4PHI3X2_MC_L5L6_L3D4),
.read_add_allprojin(AP_L5L6_L3D4_MC_L5L6_L3D4_read_add),
.allprojin(AP_L5L6_L3D4_MC_L5L6_L3D4),
.read_add_allstubin(AS_L3D4n2_MC_L5L6_L3D4_read_add),
.allstubin(AS_L3D4n2_MC_L5L6_L3D4),
.matchoutminus(MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus),
.matchoutplus(MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus),
.matchout1(MC_L5L6_L3D4_FM_L5L6_L3D4),
.valid_matchminus(MC_L5L6_L3D4_FM_L5L6_L3D4_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L3D4_FM_L5L6_L3D4_ToPlus_wr_en),
.valid_match(MC_L5L6_L3D4_FM_L5L6_L3D4_wr_en),
.start(CM_L5L6_L3D4PHI1X1_start),
.done(MC_L5L6_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b0,`PHI_L4,`Z_L4,`R_L4,`PHID_L4,`ZD_L4,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L5L6_L4,`MC_z_L5L6_L4,`MC_zfactor_OUTER) MC_L5L6_L4D3(
.number_in_match1in(CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3_number),
.read_add_match1in(CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3_read_add),
.match1in(CM_L5L6_L4D3PHI1X1_MC_L5L6_L4D3),
.number_in_match2in(CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3_number),
.read_add_match2in(CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3_read_add),
.match2in(CM_L5L6_L4D3PHI1X2_MC_L5L6_L4D3),
.number_in_match3in(CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3_number),
.read_add_match3in(CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3_read_add),
.match3in(CM_L5L6_L4D3PHI2X1_MC_L5L6_L4D3),
.number_in_match4in(CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3_number),
.read_add_match4in(CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3_read_add),
.match4in(CM_L5L6_L4D3PHI2X2_MC_L5L6_L4D3),
.number_in_match5in(CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3_number),
.read_add_match5in(CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3_read_add),
.match5in(CM_L5L6_L4D3PHI3X1_MC_L5L6_L4D3),
.number_in_match6in(CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3_number),
.read_add_match6in(CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3_read_add),
.match6in(CM_L5L6_L4D3PHI3X2_MC_L5L6_L4D3),
.number_in_match7in(CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3_number),
.read_add_match7in(CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3_read_add),
.match7in(CM_L5L6_L4D3PHI4X1_MC_L5L6_L4D3),
.number_in_match8in(CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3_number),
.read_add_match8in(CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3_read_add),
.match8in(CM_L5L6_L4D3PHI4X2_MC_L5L6_L4D3),
.read_add_allprojin(AP_L5L6_L4D3_MC_L5L6_L4D3_read_add),
.allprojin(AP_L5L6_L4D3_MC_L5L6_L4D3),
.read_add_allstubin(AS_L4D3n2_MC_L5L6_L4D3_read_add),
.allstubin(AS_L4D3n2_MC_L5L6_L4D3),
.matchoutminus(MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus),
.matchoutplus(MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus),
.matchout1(MC_L5L6_L4D3_FM_L5L6_L4D3),
.valid_matchminus(MC_L5L6_L4D3_FM_L5L6_L4D3_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L4D3_FM_L5L6_L4D3_ToPlus_wr_en),
.valid_match(MC_L5L6_L4D3_FM_L5L6_L4D3_wr_en),
.start(CM_L5L6_L4D3PHI1X1_start),
.done(MC_L5L6_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b0,`PHI_L4,`Z_L4,`R_L4,`PHID_L4,`ZD_L4,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L5L6_L4,`MC_z_L5L6_L4,`MC_zfactor_OUTER) MC_L5L6_L4D4(
.number_in_match1in(CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4_number),
.read_add_match1in(CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4_read_add),
.match1in(CM_L5L6_L4D4PHI1X1_MC_L5L6_L4D4),
.number_in_match2in(CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4_number),
.read_add_match2in(CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4_read_add),
.match2in(CM_L5L6_L4D4PHI1X2_MC_L5L6_L4D4),
.number_in_match3in(CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4_number),
.read_add_match3in(CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4_read_add),
.match3in(CM_L5L6_L4D4PHI2X1_MC_L5L6_L4D4),
.number_in_match4in(CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4_number),
.read_add_match4in(CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4_read_add),
.match4in(CM_L5L6_L4D4PHI2X2_MC_L5L6_L4D4),
.number_in_match5in(CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4_number),
.read_add_match5in(CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4_read_add),
.match5in(CM_L5L6_L4D4PHI3X1_MC_L5L6_L4D4),
.number_in_match6in(CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4_number),
.read_add_match6in(CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4_read_add),
.match6in(CM_L5L6_L4D4PHI3X2_MC_L5L6_L4D4),
.number_in_match7in(CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4_number),
.read_add_match7in(CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4_read_add),
.match7in(CM_L5L6_L4D4PHI4X1_MC_L5L6_L4D4),
.number_in_match8in(CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4_number),
.read_add_match8in(CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4_read_add),
.match8in(CM_L5L6_L4D4PHI4X2_MC_L5L6_L4D4),
.read_add_allprojin(AP_L5L6_L4D4_MC_L5L6_L4D4_read_add),
.allprojin(AP_L5L6_L4D4_MC_L5L6_L4D4),
.read_add_allstubin(AS_L4D4n3_MC_L5L6_L4D4_read_add),
.allstubin(AS_L4D4n3_MC_L5L6_L4D4),
.matchoutminus(MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus),
.matchoutplus(MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus),
.matchout1(MC_L5L6_L4D4_FM_L5L6_L4D4),
.valid_matchminus(MC_L5L6_L4D4_FM_L5L6_L4D4_ToMinus_wr_en),
.valid_matchplus(MC_L5L6_L4D4_FM_L5L6_L4D4_ToPlus_wr_en),
.valid_match(MC_L5L6_L4D4_FM_L5L6_L4D4_wr_en),
.start(CM_L5L6_L4D4PHI1X1_start),
.done(MC_L5L6_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b1,`PHI_L3,`Z_L3,`R_L3,`PHID_L3,`ZD_L3,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L1L2_L3,`MC_z_L1L2_L3,`MC_zfactor_INNER) MC_L1L2_L3D3(
.number_in_match1in(CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3_number),
.read_add_match1in(CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3_read_add),
.match1in(CM_L1L2_L3D3PHI1X1_MC_L1L2_L3D3),
.number_in_match2in(CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3_number),
.read_add_match2in(CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3_read_add),
.match2in(CM_L1L2_L3D3PHI1X2_MC_L1L2_L3D3),
.number_in_match3in(CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3_number),
.read_add_match3in(CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3_read_add),
.match3in(CM_L1L2_L3D3PHI2X1_MC_L1L2_L3D3),
.number_in_match4in(CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3_number),
.read_add_match4in(CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3_read_add),
.match4in(CM_L1L2_L3D3PHI2X2_MC_L1L2_L3D3),
.number_in_match5in(CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3_number),
.read_add_match5in(CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3_read_add),
.match5in(CM_L1L2_L3D3PHI3X1_MC_L1L2_L3D3),
.number_in_match6in(CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3_number),
.read_add_match6in(CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3_read_add),
.match6in(CM_L1L2_L3D3PHI3X2_MC_L1L2_L3D3),
.read_add_allprojin(AP_L1L2_L3D3_MC_L1L2_L3D3_read_add),
.allprojin(AP_L1L2_L3D3_MC_L1L2_L3D3),
.read_add_allstubin(AS_L3D3n4_MC_L1L2_L3D3_read_add),
.allstubin(AS_L3D3n4_MC_L1L2_L3D3),
.matchoutminus(MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus),
.matchoutplus(MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus),
.matchout1(MC_L1L2_L3D3_FM_L1L2_L3D3),
.valid_matchminus(MC_L1L2_L3D3_FM_L1L2_L3D3_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L3D3_FM_L1L2_L3D3_ToPlus_wr_en),
.valid_match(MC_L1L2_L3D3_FM_L1L2_L3D3_wr_en),
.start(CM_L1L2_L3D3PHI1X1_start),
.done(MC_L1L2_L3D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b1,`PHI_L3,`Z_L3,`R_L3,`PHID_L3,`ZD_L3,`MC_k1ABC_INNER,`MC_k2ABC_INNER,`MC_phi_L1L2_L3,`MC_z_L1L2_L3,`MC_zfactor_INNER) MC_L1L2_L3D4(
.number_in_match1in(CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4_number),
.read_add_match1in(CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4_read_add),
.match1in(CM_L1L2_L3D4PHI1X1_MC_L1L2_L3D4),
.number_in_match2in(CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4_number),
.read_add_match2in(CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4_read_add),
.match2in(CM_L1L2_L3D4PHI1X2_MC_L1L2_L3D4),
.number_in_match3in(CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4_number),
.read_add_match3in(CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4_read_add),
.match3in(CM_L1L2_L3D4PHI2X1_MC_L1L2_L3D4),
.number_in_match4in(CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4_number),
.read_add_match4in(CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4_read_add),
.match4in(CM_L1L2_L3D4PHI2X2_MC_L1L2_L3D4),
.number_in_match5in(CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4_number),
.read_add_match5in(CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4_read_add),
.match5in(CM_L1L2_L3D4PHI3X1_MC_L1L2_L3D4),
.number_in_match6in(CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4_number),
.read_add_match6in(CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4_read_add),
.match6in(CM_L1L2_L3D4PHI3X2_MC_L1L2_L3D4),
.read_add_allprojin(AP_L1L2_L3D4_MC_L1L2_L3D4_read_add),
.allprojin(AP_L1L2_L3D4_MC_L1L2_L3D4),
.read_add_allstubin(AS_L3D4n3_MC_L1L2_L3D4_read_add),
.allstubin(AS_L3D4n3_MC_L1L2_L3D4),
.matchoutminus(MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus),
.matchoutplus(MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus),
.matchout1(MC_L1L2_L3D4_FM_L1L2_L3D4),
.valid_matchminus(MC_L1L2_L3D4_FM_L1L2_L3D4_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L3D4_FM_L1L2_L3D4_ToPlus_wr_en),
.valid_match(MC_L1L2_L3D4_FM_L1L2_L3D4_wr_en),
.start(CM_L1L2_L3D4PHI1X1_start),
.done(MC_L1L2_L3D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b0,`PHI_L4,`Z_L4,`R_L4,`PHID_L4,`ZD_L4,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L4,`MC_z_L1L2_L4,`MC_zfactor_OUTER) MC_L1L2_L4D3(
.number_in_match1in(CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3_number),
.read_add_match1in(CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3_read_add),
.match1in(CM_L1L2_L4D3PHI1X1_MC_L1L2_L4D3),
.number_in_match2in(CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3_number),
.read_add_match2in(CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3_read_add),
.match2in(CM_L1L2_L4D3PHI1X2_MC_L1L2_L4D3),
.number_in_match3in(CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3_number),
.read_add_match3in(CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3_read_add),
.match3in(CM_L1L2_L4D3PHI2X1_MC_L1L2_L4D3),
.number_in_match4in(CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3_number),
.read_add_match4in(CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3_read_add),
.match4in(CM_L1L2_L4D3PHI2X2_MC_L1L2_L4D3),
.number_in_match5in(CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3_number),
.read_add_match5in(CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3_read_add),
.match5in(CM_L1L2_L4D3PHI3X1_MC_L1L2_L4D3),
.number_in_match6in(CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3_number),
.read_add_match6in(CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3_read_add),
.match6in(CM_L1L2_L4D3PHI3X2_MC_L1L2_L4D3),
.number_in_match7in(CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3_number),
.read_add_match7in(CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3_read_add),
.match7in(CM_L1L2_L4D3PHI4X1_MC_L1L2_L4D3),
.number_in_match8in(CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3_number),
.read_add_match8in(CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3_read_add),
.match8in(CM_L1L2_L4D3PHI4X2_MC_L1L2_L4D3),
.read_add_allprojin(AP_L1L2_L4D3_MC_L1L2_L4D3_read_add),
.allprojin(AP_L1L2_L4D3_MC_L1L2_L4D3),
.read_add_allstubin(AS_L4D3n3_MC_L1L2_L4D3_read_add),
.allstubin(AS_L4D3n3_MC_L1L2_L4D3),
.matchoutminus(MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus),
.matchoutplus(MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus),
.matchout1(MC_L1L2_L4D3_FM_L1L2_L4D3),
.valid_matchminus(MC_L1L2_L4D3_FM_L1L2_L4D3_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L4D3_FM_L1L2_L4D3_ToPlus_wr_en),
.valid_match(MC_L1L2_L4D3_FM_L1L2_L4D3_wr_en),
.start(CM_L1L2_L4D3PHI1X1_start),
.done(MC_L1L2_L4D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b0,`PHI_L4,`Z_L4,`R_L4,`PHID_L4,`ZD_L4,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L4,`MC_z_L1L2_L4,`MC_zfactor_OUTER) MC_L1L2_L4D4(
.number_in_match1in(CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4_number),
.read_add_match1in(CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4_read_add),
.match1in(CM_L1L2_L4D4PHI1X1_MC_L1L2_L4D4),
.number_in_match2in(CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4_number),
.read_add_match2in(CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4_read_add),
.match2in(CM_L1L2_L4D4PHI1X2_MC_L1L2_L4D4),
.number_in_match3in(CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4_number),
.read_add_match3in(CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4_read_add),
.match3in(CM_L1L2_L4D4PHI2X1_MC_L1L2_L4D4),
.number_in_match4in(CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4_number),
.read_add_match4in(CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4_read_add),
.match4in(CM_L1L2_L4D4PHI2X2_MC_L1L2_L4D4),
.number_in_match5in(CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4_number),
.read_add_match5in(CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4_read_add),
.match5in(CM_L1L2_L4D4PHI3X1_MC_L1L2_L4D4),
.number_in_match6in(CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4_number),
.read_add_match6in(CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4_read_add),
.match6in(CM_L1L2_L4D4PHI3X2_MC_L1L2_L4D4),
.number_in_match7in(CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4_number),
.read_add_match7in(CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4_read_add),
.match7in(CM_L1L2_L4D4PHI4X1_MC_L1L2_L4D4),
.number_in_match8in(CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4_number),
.read_add_match8in(CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4_read_add),
.match8in(CM_L1L2_L4D4PHI4X2_MC_L1L2_L4D4),
.read_add_allprojin(AP_L1L2_L4D4_MC_L1L2_L4D4_read_add),
.allprojin(AP_L1L2_L4D4_MC_L1L2_L4D4),
.read_add_allstubin(AS_L4D4n4_MC_L1L2_L4D4_read_add),
.allstubin(AS_L4D4n4_MC_L1L2_L4D4),
.matchoutminus(MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus),
.matchoutplus(MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus),
.matchout1(MC_L1L2_L4D4_FM_L1L2_L4D4),
.valid_matchminus(MC_L1L2_L4D4_FM_L1L2_L4D4_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L4D4_FM_L1L2_L4D4_ToPlus_wr_en),
.valid_match(MC_L1L2_L4D4_FM_L1L2_L4D4_wr_en),
.start(CM_L1L2_L4D4PHI1X1_start),
.done(MC_L1L2_L4D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b0,`PHI_L5,`Z_L5,`R_L5,`PHID_L5,`ZD_L5,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L5,`MC_z_L1L2_L5,`MC_zfactor_OUTER) MC_L1L2_L5D3(
.number_in_match1in(CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3_number),
.read_add_match1in(CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3_read_add),
.match1in(CM_L1L2_L5D3PHI1X1_MC_L1L2_L5D3),
.number_in_match2in(CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3_number),
.read_add_match2in(CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3_read_add),
.match2in(CM_L1L2_L5D3PHI1X2_MC_L1L2_L5D3),
.number_in_match3in(CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3_number),
.read_add_match3in(CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3_read_add),
.match3in(CM_L1L2_L5D3PHI2X1_MC_L1L2_L5D3),
.number_in_match4in(CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3_number),
.read_add_match4in(CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3_read_add),
.match4in(CM_L1L2_L5D3PHI2X2_MC_L1L2_L5D3),
.number_in_match5in(CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3_number),
.read_add_match5in(CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3_read_add),
.match5in(CM_L1L2_L5D3PHI3X1_MC_L1L2_L5D3),
.number_in_match6in(CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3_number),
.read_add_match6in(CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3_read_add),
.match6in(CM_L1L2_L5D3PHI3X2_MC_L1L2_L5D3),
.read_add_allprojin(AP_L1L2_L5D3_MC_L1L2_L5D3_read_add),
.allprojin(AP_L1L2_L5D3_MC_L1L2_L5D3),
.read_add_allstubin(AS_L5D3n4_MC_L1L2_L5D3_read_add),
.allstubin(AS_L5D3n4_MC_L1L2_L5D3),
.matchoutminus(MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus),
.matchoutplus(MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus),
.matchout1(MC_L1L2_L5D3_FM_L1L2_L5D3),
.valid_matchminus(MC_L1L2_L5D3_FM_L1L2_L5D3_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L5D3_FM_L1L2_L5D3_ToPlus_wr_en),
.valid_match(MC_L1L2_L5D3_FM_L1L2_L5D3_wr_en),
.start(CM_L1L2_L5D3PHI1X1_start),
.done(MC_L1L2_L5D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b0,`PHI_L5,`Z_L5,`R_L5,`PHID_L5,`ZD_L5,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L5,`MC_z_L1L2_L5,`MC_zfactor_OUTER) MC_L1L2_L5D4(
.number_in_match1in(CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4_number),
.read_add_match1in(CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4_read_add),
.match1in(CM_L1L2_L5D4PHI1X1_MC_L1L2_L5D4),
.number_in_match2in(CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4_number),
.read_add_match2in(CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4_read_add),
.match2in(CM_L1L2_L5D4PHI1X2_MC_L1L2_L5D4),
.number_in_match3in(CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4_number),
.read_add_match3in(CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4_read_add),
.match3in(CM_L1L2_L5D4PHI2X1_MC_L1L2_L5D4),
.number_in_match4in(CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4_number),
.read_add_match4in(CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4_read_add),
.match4in(CM_L1L2_L5D4PHI2X2_MC_L1L2_L5D4),
.number_in_match5in(CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4_number),
.read_add_match5in(CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4_read_add),
.match5in(CM_L1L2_L5D4PHI3X1_MC_L1L2_L5D4),
.number_in_match6in(CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4_number),
.read_add_match6in(CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4_read_add),
.match6in(CM_L1L2_L5D4PHI3X2_MC_L1L2_L5D4),
.read_add_allprojin(AP_L1L2_L5D4_MC_L1L2_L5D4_read_add),
.allprojin(AP_L1L2_L5D4_MC_L1L2_L5D4),
.read_add_allstubin(AS_L5D4n3_MC_L1L2_L5D4_read_add),
.allstubin(AS_L5D4n3_MC_L1L2_L5D4),
.matchoutminus(MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus),
.matchoutplus(MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus),
.matchout1(MC_L1L2_L5D4_FM_L1L2_L5D4),
.valid_matchminus(MC_L1L2_L5D4_FM_L1L2_L5D4_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L5D4_FM_L1L2_L5D4_ToPlus_wr_en),
.valid_match(MC_L1L2_L5D4_FM_L1L2_L5D4_wr_en),
.start(CM_L1L2_L5D4PHI1X1_start),
.done(MC_L1L2_L5D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b010,1'b0,`PHI_L6,`Z_L6,`R_L6,`PHID_L6,`ZD_L6,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L6,`MC_z_L1L2_L6,`MC_zfactor_OUTER) MC_L1L2_L6D3(
.number_in_match1in(CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3_number),
.read_add_match1in(CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3_read_add),
.match1in(CM_L1L2_L6D3PHI1X1_MC_L1L2_L6D3),
.number_in_match2in(CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3_number),
.read_add_match2in(CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3_read_add),
.match2in(CM_L1L2_L6D3PHI1X2_MC_L1L2_L6D3),
.number_in_match3in(CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3_number),
.read_add_match3in(CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3_read_add),
.match3in(CM_L1L2_L6D3PHI2X1_MC_L1L2_L6D3),
.number_in_match4in(CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3_number),
.read_add_match4in(CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3_read_add),
.match4in(CM_L1L2_L6D3PHI2X2_MC_L1L2_L6D3),
.number_in_match5in(CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3_number),
.read_add_match5in(CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3_read_add),
.match5in(CM_L1L2_L6D3PHI3X1_MC_L1L2_L6D3),
.number_in_match6in(CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3_number),
.read_add_match6in(CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3_read_add),
.match6in(CM_L1L2_L6D3PHI3X2_MC_L1L2_L6D3),
.number_in_match7in(CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3_number),
.read_add_match7in(CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3_read_add),
.match7in(CM_L1L2_L6D3PHI4X1_MC_L1L2_L6D3),
.number_in_match8in(CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3_number),
.read_add_match8in(CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3_read_add),
.match8in(CM_L1L2_L6D3PHI4X2_MC_L1L2_L6D3),
.read_add_allprojin(AP_L1L2_L6D3_MC_L1L2_L6D3_read_add),
.allprojin(AP_L1L2_L6D3_MC_L1L2_L6D3),
.read_add_allstubin(AS_L6D3n3_MC_L1L2_L6D3_read_add),
.allstubin(AS_L6D3n3_MC_L1L2_L6D3),
.matchoutminus(MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus),
.matchoutplus(MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus),
.matchout1(MC_L1L2_L6D3_FM_L1L2_L6D3),
.valid_matchminus(MC_L1L2_L6D3_FM_L1L2_L6D3_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L6D3_FM_L1L2_L6D3_ToPlus_wr_en),
.valid_match(MC_L1L2_L6D3_FM_L1L2_L6D3_wr_en),
.start(CM_L1L2_L6D3PHI1X1_start),
.done(MC_L1L2_L6D3_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchCalculator #(3'b011,1'b0,`PHI_L6,`Z_L6,`R_L6,`PHID_L6,`ZD_L6,`MC_k1ABC_OUTER,`MC_k2ABC_OUTER,`MC_phi_L1L2_L6,`MC_z_L1L2_L6,`MC_zfactor_OUTER) MC_L1L2_L6D4(
.number_in_match1in(CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4_number),
.read_add_match1in(CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4_read_add),
.match1in(CM_L1L2_L6D4PHI1X1_MC_L1L2_L6D4),
.number_in_match2in(CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4_number),
.read_add_match2in(CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4_read_add),
.match2in(CM_L1L2_L6D4PHI1X2_MC_L1L2_L6D4),
.number_in_match3in(CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4_number),
.read_add_match3in(CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4_read_add),
.match3in(CM_L1L2_L6D4PHI2X1_MC_L1L2_L6D4),
.number_in_match4in(CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4_number),
.read_add_match4in(CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4_read_add),
.match4in(CM_L1L2_L6D4PHI2X2_MC_L1L2_L6D4),
.number_in_match5in(CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4_number),
.read_add_match5in(CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4_read_add),
.match5in(CM_L1L2_L6D4PHI3X1_MC_L1L2_L6D4),
.number_in_match6in(CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4_number),
.read_add_match6in(CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4_read_add),
.match6in(CM_L1L2_L6D4PHI3X2_MC_L1L2_L6D4),
.number_in_match7in(CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4_number),
.read_add_match7in(CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4_read_add),
.match7in(CM_L1L2_L6D4PHI4X1_MC_L1L2_L6D4),
.number_in_match8in(CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4_number),
.read_add_match8in(CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4_read_add),
.match8in(CM_L1L2_L6D4PHI4X2_MC_L1L2_L6D4),
.read_add_allprojin(AP_L1L2_L6D4_MC_L1L2_L6D4_read_add),
.allprojin(AP_L1L2_L6D4_MC_L1L2_L6D4),
.read_add_allstubin(AS_L6D4n4_MC_L1L2_L6D4_read_add),
.allstubin(AS_L6D4n4_MC_L1L2_L6D4),
.matchoutminus(MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus),
.matchoutplus(MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus),
.matchout1(MC_L1L2_L6D4_FM_L1L2_L6D4),
.valid_matchminus(MC_L1L2_L6D4_FM_L1L2_L6D4_ToMinus_wr_en),
.valid_matchplus(MC_L1L2_L6D4_FM_L1L2_L6D4_ToPlus_wr_en),
.valid_match(MC_L1L2_L6D4_FM_L1L2_L6D4_wr_en),
.start(CM_L1L2_L6D4PHI1X1_start),
.done(MC_L1L2_L6D4_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchTransceiver #("Layer") MT_Layr_Minus(
.number_in1(FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_number),
.read_add1(FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_read_add),
.read_en1(FM_L1L2_L3D3_ToMinus_MT_Layr_Minus_read_en),
.matchin1(FM_L1L2_L3D3_ToMinus_MT_Layr_Minus),
.number_in2(FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_number),
.read_add2(FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_read_add),
.read_en2(FM_L1L2_L4D3_ToMinus_MT_Layr_Minus_read_en),
.matchin2(FM_L1L2_L4D3_ToMinus_MT_Layr_Minus),
.number_in3(FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_number),
.read_add3(FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_read_add),
.read_en3(FM_L1L2_L5D3_ToMinus_MT_Layr_Minus_read_en),
.matchin3(FM_L1L2_L5D3_ToMinus_MT_Layr_Minus),
.number_in4(FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_number),
.read_add4(FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_read_add),
.read_en4(FM_L1L2_L6D3_ToMinus_MT_Layr_Minus_read_en),
.matchin4(FM_L1L2_L6D3_ToMinus_MT_Layr_Minus),
.number_in5(FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_number),
.read_add5(FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_read_add),
.read_en5(FM_L3L4_L1D3_ToMinus_MT_Layr_Minus_read_en),
.matchin5(FM_L3L4_L1D3_ToMinus_MT_Layr_Minus),
.number_in6(FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_number),
.read_add6(FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_read_add),
.read_en6(FM_L3L4_L2D3_ToMinus_MT_Layr_Minus_read_en),
.matchin6(FM_L3L4_L2D3_ToMinus_MT_Layr_Minus),
.number_in7(FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_number),
.read_add7(FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_read_add),
.read_en7(FM_L3L4_L5D3_ToMinus_MT_Layr_Minus_read_en),
.matchin7(FM_L3L4_L5D3_ToMinus_MT_Layr_Minus),
.number_in8(FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_number),
.read_add8(FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_read_add),
.read_en8(FM_L3L4_L6D3_ToMinus_MT_Layr_Minus_read_en),
.matchin8(FM_L3L4_L6D3_ToMinus_MT_Layr_Minus),
.number_in9(FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_number),
.read_add9(FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_read_add),
.read_en9(FM_L5L6_L1D3_ToMinus_MT_Layr_Minus_read_en),
.matchin9(FM_L5L6_L1D3_ToMinus_MT_Layr_Minus),
.number_in10(FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_number),
.read_add10(FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_read_add),
.read_en10(FM_L5L6_L2D3_ToMinus_MT_Layr_Minus_read_en),
.matchin10(FM_L5L6_L2D3_ToMinus_MT_Layr_Minus),
.number_in11(FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_number),
.read_add11(FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_read_add),
.read_en11(FM_L5L6_L3D3_ToMinus_MT_Layr_Minus_read_en),
.matchin11(FM_L5L6_L3D3_ToMinus_MT_Layr_Minus),
.number_in12(FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_number),
.read_add12(FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_read_add),
.read_en12(FM_L5L6_L4D3_ToMinus_MT_Layr_Minus_read_en),
.matchin12(FM_L5L6_L4D3_ToMinus_MT_Layr_Minus),
.number_in13(FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_number),
.read_add13(FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_read_add),
.read_en13(FM_L1L2_L3D4_ToMinus_MT_Layr_Minus_read_en),
.matchin13(FM_L1L2_L3D4_ToMinus_MT_Layr_Minus),
.number_in14(FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_number),
.read_add14(FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_read_add),
.read_en14(FM_L1L2_L4D4_ToMinus_MT_Layr_Minus_read_en),
.matchin14(FM_L1L2_L4D4_ToMinus_MT_Layr_Minus),
.number_in15(FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_number),
.read_add15(FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_read_add),
.read_en15(FM_L1L2_L5D4_ToMinus_MT_Layr_Minus_read_en),
.matchin15(FM_L1L2_L5D4_ToMinus_MT_Layr_Minus),
.number_in16(FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_number),
.read_add16(FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_read_add),
.read_en16(FM_L1L2_L6D4_ToMinus_MT_Layr_Minus_read_en),
.matchin16(FM_L1L2_L6D4_ToMinus_MT_Layr_Minus),
.number_in17(FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_number),
.read_add17(FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_read_add),
.read_en17(FM_L3L4_L1D4_ToMinus_MT_Layr_Minus_read_en),
.matchin17(FM_L3L4_L1D4_ToMinus_MT_Layr_Minus),
.number_in18(FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_number),
.read_add18(FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_read_add),
.read_en18(FM_L3L4_L2D4_ToMinus_MT_Layr_Minus_read_en),
.matchin18(FM_L3L4_L2D4_ToMinus_MT_Layr_Minus),
.number_in19(FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_number),
.read_add19(FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_read_add),
.read_en19(FM_L3L4_L5D4_ToMinus_MT_Layr_Minus_read_en),
.matchin19(FM_L3L4_L5D4_ToMinus_MT_Layr_Minus),
.number_in20(FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_number),
.read_add20(FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_read_add),
.read_en20(FM_L3L4_L6D4_ToMinus_MT_Layr_Minus_read_en),
.matchin20(FM_L3L4_L6D4_ToMinus_MT_Layr_Minus),
.number_in21(FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_number),
.read_add21(FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_read_add),
.read_en21(FM_L5L6_L1D4_ToMinus_MT_Layr_Minus_read_en),
.matchin21(FM_L5L6_L1D4_ToMinus_MT_Layr_Minus),
.number_in22(FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_number),
.read_add22(FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_read_add),
.read_en22(FM_L5L6_L2D4_ToMinus_MT_Layr_Minus_read_en),
.matchin22(FM_L5L6_L2D4_ToMinus_MT_Layr_Minus),
.number_in23(FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_number),
.read_add23(FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_read_add),
.read_en23(FM_L5L6_L3D4_ToMinus_MT_Layr_Minus_read_en),
.matchin23(FM_L5L6_L3D4_ToMinus_MT_Layr_Minus),
.number_in24(FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_number),
.read_add24(FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_read_add),
.read_en24(FM_L5L6_L4D4_ToMinus_MT_Layr_Minus_read_en),
.matchin24(FM_L5L6_L4D4_ToMinus_MT_Layr_Minus),
.valid_incomming_match_data_stream(MT_Layr_Minus_From_DataStream_en),
.incomming_match_data_stream(MT_Layr_Minus_From_DataStream),
.matchout1(MT_Layr_Minus_FM_L1L2_L3_FromMinus),
.matchout2(MT_Layr_Minus_FM_L1L2_L4_FromMinus),
.matchout3(MT_Layr_Minus_FM_L1L2_L5_FromMinus),
.matchout4(MT_Layr_Minus_FM_L1L2_L6_FromMinus),
.matchout5(MT_Layr_Minus_FM_L3L4_L1_FromMinus),
.matchout6(MT_Layr_Minus_FM_L3L4_L2_FromMinus),
.matchout7(MT_Layr_Minus_FM_L3L4_L5_FromMinus),
.matchout8(MT_Layr_Minus_FM_L3L4_L6_FromMinus),
.matchout9(MT_Layr_Minus_FM_L5L6_L1_FromMinus),
.matchout10(MT_Layr_Minus_FM_L5L6_L2_FromMinus),
.matchout11(MT_Layr_Minus_FM_L5L6_L3_FromMinus),
.matchout12(MT_Layr_Minus_FM_L5L6_L4_FromMinus),
.valid_matchout1(MT_Layr_Minus_FM_L1L2_L3_FromMinus_wr_en),
.valid_matchout2(MT_Layr_Minus_FM_L1L2_L4_FromMinus_wr_en),
.valid_matchout3(MT_Layr_Minus_FM_L1L2_L5_FromMinus_wr_en),
.valid_matchout4(MT_Layr_Minus_FM_L1L2_L6_FromMinus_wr_en),
.valid_matchout5(MT_Layr_Minus_FM_L3L4_L1_FromMinus_wr_en),
.valid_matchout6(MT_Layr_Minus_FM_L3L4_L2_FromMinus_wr_en),
.valid_matchout7(MT_Layr_Minus_FM_L3L4_L5_FromMinus_wr_en),
.valid_matchout8(MT_Layr_Minus_FM_L3L4_L6_FromMinus_wr_en),
.valid_matchout9(MT_Layr_Minus_FM_L5L6_L1_FromMinus_wr_en),
.valid_matchout10(MT_Layr_Minus_FM_L5L6_L2_FromMinus_wr_en),
.valid_matchout11(MT_Layr_Minus_FM_L5L6_L3_FromMinus_wr_en),
.valid_matchout12(MT_Layr_Minus_FM_L5L6_L4_FromMinus_wr_en),
.valid_match_data_stream(MT_Layr_Minus_To_DataStream_en),
.match_data_stream(MT_Layr_Minus_To_DataStream),
.start(FM_L1L2_L3D3_ToMinus_start),
.done(MT_Layr_Minus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

MatchTransceiver #("Layer") MT_Layr_Plus(
.number_in1(FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_number),
.read_add1(FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_read_add),
.read_en1(FM_L1L2_L3D3_ToPlus_MT_Layr_Plus_read_en),
.matchin1(FM_L1L2_L3D3_ToPlus_MT_Layr_Plus),
.number_in2(FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_number),
.read_add2(FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_read_add),
.read_en2(FM_L1L2_L4D3_ToPlus_MT_Layr_Plus_read_en),
.matchin2(FM_L1L2_L4D3_ToPlus_MT_Layr_Plus),
.number_in3(FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_number),
.read_add3(FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_read_add),
.read_en3(FM_L1L2_L5D3_ToPlus_MT_Layr_Plus_read_en),
.matchin3(FM_L1L2_L5D3_ToPlus_MT_Layr_Plus),
.number_in4(FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_number),
.read_add4(FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_read_add),
.read_en4(FM_L1L2_L6D3_ToPlus_MT_Layr_Plus_read_en),
.matchin4(FM_L1L2_L6D3_ToPlus_MT_Layr_Plus),
.number_in5(FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_number),
.read_add5(FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_read_add),
.read_en5(FM_L3L4_L1D3_ToPlus_MT_Layr_Plus_read_en),
.matchin5(FM_L3L4_L1D3_ToPlus_MT_Layr_Plus),
.number_in6(FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_number),
.read_add6(FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_read_add),
.read_en6(FM_L3L4_L2D3_ToPlus_MT_Layr_Plus_read_en),
.matchin6(FM_L3L4_L2D3_ToPlus_MT_Layr_Plus),
.number_in7(FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_number),
.read_add7(FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_read_add),
.read_en7(FM_L3L4_L5D3_ToPlus_MT_Layr_Plus_read_en),
.matchin7(FM_L3L4_L5D3_ToPlus_MT_Layr_Plus),
.number_in8(FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_number),
.read_add8(FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_read_add),
.read_en8(FM_L3L4_L6D3_ToPlus_MT_Layr_Plus_read_en),
.matchin8(FM_L3L4_L6D3_ToPlus_MT_Layr_Plus),
.number_in9(FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_number),
.read_add9(FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_read_add),
.read_en9(FM_L5L6_L1D3_ToPlus_MT_Layr_Plus_read_en),
.matchin9(FM_L5L6_L1D3_ToPlus_MT_Layr_Plus),
.number_in10(FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_number),
.read_add10(FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_read_add),
.read_en10(FM_L5L6_L2D3_ToPlus_MT_Layr_Plus_read_en),
.matchin10(FM_L5L6_L2D3_ToPlus_MT_Layr_Plus),
.number_in11(FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_number),
.read_add11(FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_read_add),
.read_en11(FM_L5L6_L3D3_ToPlus_MT_Layr_Plus_read_en),
.matchin11(FM_L5L6_L3D3_ToPlus_MT_Layr_Plus),
.number_in12(FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_number),
.read_add12(FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_read_add),
.read_en12(FM_L5L6_L4D3_ToPlus_MT_Layr_Plus_read_en),
.matchin12(FM_L5L6_L4D3_ToPlus_MT_Layr_Plus),
.number_in13(FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_number),
.read_add13(FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_read_add),
.read_en13(FM_L1L2_L3D4_ToPlus_MT_Layr_Plus_read_en),
.matchin13(FM_L1L2_L3D4_ToPlus_MT_Layr_Plus),
.number_in14(FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_number),
.read_add14(FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_read_add),
.read_en14(FM_L1L2_L4D4_ToPlus_MT_Layr_Plus_read_en),
.matchin14(FM_L1L2_L4D4_ToPlus_MT_Layr_Plus),
.number_in15(FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_number),
.read_add15(FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_read_add),
.read_en15(FM_L1L2_L5D4_ToPlus_MT_Layr_Plus_read_en),
.matchin15(FM_L1L2_L5D4_ToPlus_MT_Layr_Plus),
.number_in16(FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_number),
.read_add16(FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_read_add),
.read_en16(FM_L1L2_L6D4_ToPlus_MT_Layr_Plus_read_en),
.matchin16(FM_L1L2_L6D4_ToPlus_MT_Layr_Plus),
.number_in17(FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_number),
.read_add17(FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_read_add),
.read_en17(FM_L3L4_L1D4_ToPlus_MT_Layr_Plus_read_en),
.matchin17(FM_L3L4_L1D4_ToPlus_MT_Layr_Plus),
.number_in18(FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_number),
.read_add18(FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_read_add),
.read_en18(FM_L3L4_L2D4_ToPlus_MT_Layr_Plus_read_en),
.matchin18(FM_L3L4_L2D4_ToPlus_MT_Layr_Plus),
.number_in19(FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_number),
.read_add19(FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_read_add),
.read_en19(FM_L3L4_L5D4_ToPlus_MT_Layr_Plus_read_en),
.matchin19(FM_L3L4_L5D4_ToPlus_MT_Layr_Plus),
.number_in20(FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_number),
.read_add20(FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_read_add),
.read_en20(FM_L3L4_L6D4_ToPlus_MT_Layr_Plus_read_en),
.matchin20(FM_L3L4_L6D4_ToPlus_MT_Layr_Plus),
.number_in21(FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_number),
.read_add21(FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_read_add),
.read_en21(FM_L5L6_L1D4_ToPlus_MT_Layr_Plus_read_en),
.matchin21(FM_L5L6_L1D4_ToPlus_MT_Layr_Plus),
.number_in22(FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_number),
.read_add22(FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_read_add),
.read_en22(FM_L5L6_L2D4_ToPlus_MT_Layr_Plus_read_en),
.matchin22(FM_L5L6_L2D4_ToPlus_MT_Layr_Plus),
.number_in23(FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_number),
.read_add23(FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_read_add),
.read_en23(FM_L5L6_L3D4_ToPlus_MT_Layr_Plus_read_en),
.matchin23(FM_L5L6_L3D4_ToPlus_MT_Layr_Plus),
.number_in24(FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_number),
.read_add24(FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_read_add),
.read_en24(FM_L5L6_L4D4_ToPlus_MT_Layr_Plus_read_en),
.matchin24(FM_L5L6_L4D4_ToPlus_MT_Layr_Plus),
.valid_incomming_match_data_stream(MT_Layr_Plus_From_DataStream_en),
.incomming_match_data_stream(MT_Layr_Plus_From_DataStream),
.matchout1(MT_Layr_Plus_FM_L1L2_L3_FromPlus),
.matchout2(MT_Layr_Plus_FM_L1L2_L4_FromPlus),
.matchout3(MT_Layr_Plus_FM_L1L2_L5_FromPlus),
.matchout4(MT_Layr_Plus_FM_L1L2_L6_FromPlus),
.matchout5(MT_Layr_Plus_FM_L3L4_L1_FromPlus),
.matchout6(MT_Layr_Plus_FM_L3L4_L2_FromPlus),
.matchout7(MT_Layr_Plus_FM_L3L4_L5_FromPlus),
.matchout8(MT_Layr_Plus_FM_L3L4_L6_FromPlus),
.matchout9(MT_Layr_Plus_FM_L5L6_L1_FromPlus),
.matchout10(MT_Layr_Plus_FM_L5L6_L2_FromPlus),
.matchout11(MT_Layr_Plus_FM_L5L6_L3_FromPlus),
.matchout12(MT_Layr_Plus_FM_L5L6_L4_FromPlus),
.valid_matchout1(MT_Layr_Plus_FM_L1L2_L3_FromPlus_wr_en),
.valid_matchout2(MT_Layr_Plus_FM_L1L2_L4_FromPlus_wr_en),
.valid_matchout3(MT_Layr_Plus_FM_L1L2_L5_FromPlus_wr_en),
.valid_matchout4(MT_Layr_Plus_FM_L1L2_L6_FromPlus_wr_en),
.valid_matchout5(MT_Layr_Plus_FM_L3L4_L1_FromPlus_wr_en),
.valid_matchout6(MT_Layr_Plus_FM_L3L4_L2_FromPlus_wr_en),
.valid_matchout7(MT_Layr_Plus_FM_L3L4_L5_FromPlus_wr_en),
.valid_matchout8(MT_Layr_Plus_FM_L3L4_L6_FromPlus_wr_en),
.valid_matchout9(MT_Layr_Plus_FM_L5L6_L1_FromPlus_wr_en),
.valid_matchout10(MT_Layr_Plus_FM_L5L6_L2_FromPlus_wr_en),
.valid_matchout11(MT_Layr_Plus_FM_L5L6_L3_FromPlus_wr_en),
.valid_matchout12(MT_Layr_Plus_FM_L5L6_L4_FromPlus_wr_en),
.valid_match_data_stream(MT_Layr_Plus_To_DataStream_en),
.match_data_stream(MT_Layr_Plus_To_DataStream),
.start(FM_L1L2_L3D3_ToPlus_start),
.done(MT_Layr_Plus_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

FitTrack #("L1L2") FT_L1L2(
.number1in1(FM_L1L2_L3D3_FT_L1L2_number),
.read_add1in1(FM_L1L2_L3D3_FT_L1L2_read_add),
.read_en1in1(FM_L1L2_L3D3_FT_L1L2_read_en),
.fullmatch1in1(FM_L1L2_L3D3_FT_L1L2),
.number1in2(FM_L1L2_L3D4_FT_L1L2_number),
.read_add1in2(FM_L1L2_L3D4_FT_L1L2_read_add),
.read_en1in2(FM_L1L2_L3D4_FT_L1L2_read_en),
.fullmatch1in2(FM_L1L2_L3D4_FT_L1L2),
.number2in1(FM_L1L2_L4D3_FT_L1L2_number),
.read_add2in1(FM_L1L2_L4D3_FT_L1L2_read_add),
.read_en2in1(FM_L1L2_L4D3_FT_L1L2_read_en),
.fullmatch2in1(FM_L1L2_L4D3_FT_L1L2),
.number2in2(FM_L1L2_L4D4_FT_L1L2_number),
.read_add2in2(FM_L1L2_L4D4_FT_L1L2_read_add),
.read_en2in2(FM_L1L2_L4D4_FT_L1L2_read_en),
.fullmatch2in2(FM_L1L2_L4D4_FT_L1L2),
.number3in1(FM_L1L2_L5D3_FT_L1L2_number),
.read_add3in1(FM_L1L2_L5D3_FT_L1L2_read_add),
.read_en3in1(FM_L1L2_L5D3_FT_L1L2_read_en),
.fullmatch3in1(FM_L1L2_L5D3_FT_L1L2),
.number3in2(FM_L1L2_L5D4_FT_L1L2_number),
.read_add3in2(FM_L1L2_L5D4_FT_L1L2_read_add),
.read_en3in2(FM_L1L2_L5D4_FT_L1L2_read_en),
.fullmatch3in2(FM_L1L2_L5D4_FT_L1L2),
.number4in1(FM_L1L2_L6D3_FT_L1L2_number),
.read_add4in1(FM_L1L2_L6D3_FT_L1L2_read_add),
.read_en4in1(FM_L1L2_L6D3_FT_L1L2_read_en),
.fullmatch4in1(FM_L1L2_L6D3_FT_L1L2),
.number4in2(FM_L1L2_L6D4_FT_L1L2_number),
.read_add4in2(FM_L1L2_L6D4_FT_L1L2_read_add),
.read_en4in2(FM_L1L2_L6D4_FT_L1L2_read_en),
.fullmatch4in2(FM_L1L2_L6D4_FT_L1L2),
.read_add_pars1(TPAR_L1D3L2D3_FT_L1L2_read_add),
.tpar1in(TPAR_L1D3L2D3_FT_L1L2),
.read_add_pars2(TPAR_L1D3L2D4_FT_L1L2_read_add),
.tpar2in(TPAR_L1D3L2D4_FT_L1L2),
.read_add_pars3(TPAR_L1D4L2D4_FT_L1L2_read_add),
.tpar3in(TPAR_L1D4L2D4_FT_L1L2),
.number1in3(FM_L1L2_L3_FromPlus_FT_L1L2_number),
.read_add1in3(FM_L1L2_L3_FromPlus_FT_L1L2_read_add),
.read_en1in3(FM_L1L2_L3_FromPlus_FT_L1L2_read_en),
.fullmatch1in3(FM_L1L2_L3_FromPlus_FT_L1L2),
.number2in3(FM_L1L2_L4_FromPlus_FT_L1L2_number),
.read_add2in3(FM_L1L2_L4_FromPlus_FT_L1L2_read_add),
.read_en2in3(FM_L1L2_L4_FromPlus_FT_L1L2_read_en),
.fullmatch2in3(FM_L1L2_L4_FromPlus_FT_L1L2),
.number3in3(FM_L1L2_L5_FromPlus_FT_L1L2_number),
.read_add3in3(FM_L1L2_L5_FromPlus_FT_L1L2_read_add),
.read_en3in3(FM_L1L2_L5_FromPlus_FT_L1L2_read_en),
.fullmatch3in3(FM_L1L2_L5_FromPlus_FT_L1L2),
.number4in3(FM_L1L2_L6_FromPlus_FT_L1L2_number),
.read_add4in3(FM_L1L2_L6_FromPlus_FT_L1L2_read_add),
.read_en4in3(FM_L1L2_L6_FromPlus_FT_L1L2_read_en),
.fullmatch4in3(FM_L1L2_L6_FromPlus_FT_L1L2),
.number1in4(FM_L1L2_L3_FromMinus_FT_L1L2_number),
.read_add1in4(FM_L1L2_L3_FromMinus_FT_L1L2_read_add),
.read_en1in4(FM_L1L2_L3_FromMinus_FT_L1L2_read_en),
.fullmatch1in4(FM_L1L2_L3_FromMinus_FT_L1L2),
.number2in4(FM_L1L2_L4_FromMinus_FT_L1L2_number),
.read_add2in4(FM_L1L2_L4_FromMinus_FT_L1L2_read_add),
.read_en2in4(FM_L1L2_L4_FromMinus_FT_L1L2_read_en),
.fullmatch2in4(FM_L1L2_L4_FromMinus_FT_L1L2),
.number3in4(FM_L1L2_L5_FromMinus_FT_L1L2_number),
.read_add3in4(FM_L1L2_L5_FromMinus_FT_L1L2_read_add),
.read_en3in4(FM_L1L2_L5_FromMinus_FT_L1L2_read_en),
.fullmatch3in4(FM_L1L2_L5_FromMinus_FT_L1L2),
.number4in4(FM_L1L2_L6_FromMinus_FT_L1L2_number),
.read_add4in4(FM_L1L2_L6_FromMinus_FT_L1L2_read_add),
.read_en4in4(FM_L1L2_L6_FromMinus_FT_L1L2_read_en),
.fullmatch4in4(FM_L1L2_L6_FromMinus_FT_L1L2),
.trackout(FT_L1L2_TF_L1L2),
.valid_fit(FT_L1L2_TF_L1L2_wr_en),
.start(FM_L1L2_L6_FromMinus_start),
.done(FT_L1L2_start),
.clk(clk),
.clk_new(clk_new),		  //MT			   
.reset(reset),
.en_proc(en_proc)
);

FitTrack #("L3L4") FT_L3L4(
.number1in1(FM_L3L4_L1D3_FT_L3L4_number),
.read_add1in1(FM_L3L4_L1D3_FT_L3L4_read_add),
.read_en1in1(FM_L3L4_L1D3_FT_L3L4_read_en),
.fullmatch1in1(FM_L3L4_L1D3_FT_L3L4),
.number1in2(FM_L3L4_L1D4_FT_L3L4_number),
.read_add1in2(FM_L3L4_L1D4_FT_L3L4_read_add),
.read_en1in2(FM_L3L4_L1D4_FT_L3L4_read_en),
.fullmatch1in2(FM_L3L4_L1D4_FT_L3L4),
.number2in1(FM_L3L4_L2D3_FT_L3L4_number),
.read_add2in1(FM_L3L4_L2D3_FT_L3L4_read_add),
.read_en2in1(FM_L3L4_L2D3_FT_L3L4_read_en),
.fullmatch2in1(FM_L3L4_L2D3_FT_L3L4),
.number2in2(FM_L3L4_L2D4_FT_L3L4_number),
.read_add2in2(FM_L3L4_L2D4_FT_L3L4_read_add),
.read_en2in2(FM_L3L4_L2D4_FT_L3L4_read_en),
.fullmatch2in2(FM_L3L4_L2D4_FT_L3L4),
.number3in1(FM_L3L4_L5D3_FT_L3L4_number),
.read_add3in1(FM_L3L4_L5D3_FT_L3L4_read_add),
.read_en3in1(FM_L3L4_L5D3_FT_L3L4_read_en),
.fullmatch3in1(FM_L3L4_L5D3_FT_L3L4),
.number3in2(FM_L3L4_L5D4_FT_L3L4_number),
.read_add3in2(FM_L3L4_L5D4_FT_L3L4_read_add),
.read_en3in2(FM_L3L4_L5D4_FT_L3L4_read_en),
.fullmatch3in2(FM_L3L4_L5D4_FT_L3L4),
.number4in1(FM_L3L4_L6D3_FT_L3L4_number),
.read_add4in1(FM_L3L4_L6D3_FT_L3L4_read_add),
.read_en4in1(FM_L3L4_L6D3_FT_L3L4_read_en),
.fullmatch4in1(FM_L3L4_L6D3_FT_L3L4),
.number4in2(FM_L3L4_L6D4_FT_L3L4_number),
.read_add4in2(FM_L3L4_L6D4_FT_L3L4_read_add),
.read_en4in2(FM_L3L4_L6D4_FT_L3L4_read_en),
.fullmatch4in2(FM_L3L4_L6D4_FT_L3L4),
.number1in3(FM_L3L4_L1_FromMinus_FT_L3L4_number),
.read_add1in3(FM_L3L4_L1_FromMinus_FT_L3L4_read_add),
.read_en1in3(FM_L3L4_L1_FromMinus_FT_L3L4_read_en),
.fullmatch1in3(FM_L3L4_L1_FromMinus_FT_L3L4),
.number2in3(FM_L3L4_L2_FromMinus_FT_L3L4_number),
.read_add2in3(FM_L3L4_L2_FromMinus_FT_L3L4_read_add),
.read_en2in3(FM_L3L4_L2_FromMinus_FT_L3L4_read_en),
.fullmatch2in3(FM_L3L4_L2_FromMinus_FT_L3L4),
.number3in3(FM_L3L4_L5_FromMinus_FT_L3L4_number),
.read_add3in3(FM_L3L4_L5_FromMinus_FT_L3L4_read_add),
.read_en3in3(FM_L3L4_L5_FromMinus_FT_L3L4_read_en),
.fullmatch3in3(FM_L3L4_L5_FromMinus_FT_L3L4),
.number4in3(FM_L3L4_L6_FromMinus_FT_L3L4_number),
.read_add4in3(FM_L3L4_L6_FromMinus_FT_L3L4_read_add),
.read_en4in3(FM_L3L4_L6_FromMinus_FT_L3L4_read_en),
.fullmatch4in3(FM_L3L4_L6_FromMinus_FT_L3L4),
.number1in4(FM_L3L4_L1_FromPlus_FT_L3L4_number),
.read_add1in4(FM_L3L4_L1_FromPlus_FT_L3L4_read_add),
.read_en1in4(FM_L3L4_L1_FromPlus_FT_L3L4_read_en),
.fullmatch1in4(FM_L3L4_L1_FromPlus_FT_L3L4),
.number2in4(FM_L3L4_L2_FromPlus_FT_L3L4_number),
.read_add2in4(FM_L3L4_L2_FromPlus_FT_L3L4_read_add),
.read_en2in4(FM_L3L4_L2_FromPlus_FT_L3L4_read_en),
.fullmatch2in4(FM_L3L4_L2_FromPlus_FT_L3L4),
.number3in4(FM_L3L4_L5_FromPlus_FT_L3L4_number),
.read_add3in4(FM_L3L4_L5_FromPlus_FT_L3L4_read_add),
.read_en3in4(FM_L3L4_L5_FromPlus_FT_L3L4_read_en),
.fullmatch3in4(FM_L3L4_L5_FromPlus_FT_L3L4),
.number4in4(FM_L3L4_L6_FromPlus_FT_L3L4_number),
.read_add4in4(FM_L3L4_L6_FromPlus_FT_L3L4_read_add),
.read_en4in4(FM_L3L4_L6_FromPlus_FT_L3L4_read_en),
.fullmatch4in4(FM_L3L4_L6_FromPlus_FT_L3L4),
.read_add_pars1(TPAR_L3D3L4D3_FT_L3L4_read_add),
.tpar1in(TPAR_L3D3L4D3_FT_L3L4),
.read_add_pars2(TPAR_L3D3L4D4_FT_L3L4_read_add),
.tpar2in(TPAR_L3D3L4D4_FT_L3L4),
.read_add_pars3(TPAR_L3D4L4D4_FT_L3L4_read_add),
.tpar3in(TPAR_L3D4L4D4_FT_L3L4),
.trackout(FT_L3L4_TF_L3L4),
.valid_fit(FT_L3L4_TF_L3L4_wr_en),
.start(FM_L3L4_L6_FromPlus_start),
.done(FT_L3L4_start),
.clk(clk),
.clk_new(clk_new),		  //MT			   
.reset(reset),
.en_proc(en_proc)
);

FitTrack #("L5L6") FT_L5L6(
.number1in1(FM_L5L6_L1D3_FT_L5L6_number),
.read_add1in1(FM_L5L6_L1D3_FT_L5L6_read_add),
.read_en1in1(FM_L5L6_L1D3_FT_L5L6_read_en),
.fullmatch1in1(FM_L5L6_L1D3_FT_L5L6),
.number1in2(FM_L5L6_L1D4_FT_L5L6_number),
.read_add1in2(FM_L5L6_L1D4_FT_L5L6_read_add),
.read_en1in2(FM_L5L6_L1D4_FT_L5L6_read_en),
.fullmatch1in2(FM_L5L6_L1D4_FT_L5L6),
.number2in1(FM_L5L6_L2D3_FT_L5L6_number),
.read_add2in1(FM_L5L6_L2D3_FT_L5L6_read_add),
.read_en2in1(FM_L5L6_L2D3_FT_L5L6_read_en),
.fullmatch2in1(FM_L5L6_L2D3_FT_L5L6),
.number2in2(FM_L5L6_L2D4_FT_L5L6_number),
.read_add2in2(FM_L5L6_L2D4_FT_L5L6_read_add),
.read_en2in2(FM_L5L6_L2D4_FT_L5L6_read_en),
.fullmatch2in2(FM_L5L6_L2D4_FT_L5L6),
.number3in1(FM_L5L6_L3D3_FT_L5L6_number),
.read_add3in1(FM_L5L6_L3D3_FT_L5L6_read_add),
.read_en3in1(FM_L5L6_L3D3_FT_L5L6_read_en),
.fullmatch3in1(FM_L5L6_L3D3_FT_L5L6),
.number3in2(FM_L5L6_L3D4_FT_L5L6_number),
.read_add3in2(FM_L5L6_L3D4_FT_L5L6_read_add),
.read_en3in2(FM_L5L6_L3D4_FT_L5L6_read_en),
.fullmatch3in2(FM_L5L6_L3D4_FT_L5L6),
.number4in1(FM_L5L6_L4D3_FT_L5L6_number),
.read_add4in1(FM_L5L6_L4D3_FT_L5L6_read_add),
.read_en4in1(FM_L5L6_L4D3_FT_L5L6_read_en),
.fullmatch4in1(FM_L5L6_L4D3_FT_L5L6),
.number4in2(FM_L5L6_L4D4_FT_L5L6_number),
.read_add4in2(FM_L5L6_L4D4_FT_L5L6_read_add),
.read_en4in2(FM_L5L6_L4D4_FT_L5L6_read_en),
.fullmatch4in2(FM_L5L6_L4D4_FT_L5L6),
.read_add_pars1(TPAR_L5D3L6D3_FT_L5L6_read_add),
.tpar1in(TPAR_L5D3L6D3_FT_L5L6),
.read_add_pars2(TPAR_L5D3L6D4_FT_L5L6_read_add),
.tpar2in(TPAR_L5D3L6D4_FT_L5L6),
.read_add_pars3(TPAR_L5D4L6D4_FT_L5L6_read_add),
.tpar3in(TPAR_L5D4L6D4_FT_L5L6),
.number1in3(FM_L5L6_L1_FromPlus_FT_L5L6_number),
.read_add1in3(FM_L5L6_L1_FromPlus_FT_L5L6_read_add),
.read_en1in3(FM_L5L6_L1_FromPlus_FT_L5L6_read_en),
.fullmatch1in3(FM_L5L6_L1_FromPlus_FT_L5L6),
.number2in3(FM_L5L6_L2_FromPlus_FT_L5L6_number),
.read_add2in3(FM_L5L6_L2_FromPlus_FT_L5L6_read_add),
.read_en2in3(FM_L5L6_L2_FromPlus_FT_L5L6_read_en),
.fullmatch2in3(FM_L5L6_L2_FromPlus_FT_L5L6),
.number3in3(FM_L5L6_L3_FromPlus_FT_L5L6_number),
.read_add3in3(FM_L5L6_L3_FromPlus_FT_L5L6_read_add),
.read_en3in3(FM_L5L6_L3_FromPlus_FT_L5L6_read_en),
.fullmatch3in3(FM_L5L6_L3_FromPlus_FT_L5L6),
.number4in3(FM_L5L6_L4_FromPlus_FT_L5L6_number),
.read_add4in3(FM_L5L6_L4_FromPlus_FT_L5L6_read_add),
.read_en4in3(FM_L5L6_L4_FromPlus_FT_L5L6_read_en),
.fullmatch4in3(FM_L5L6_L4_FromPlus_FT_L5L6),
.number1in4(FM_L5L6_L1_FromMinus_FT_L5L6_number),
.read_add1in4(FM_L5L6_L1_FromMinus_FT_L5L6_read_add),
.read_en1in4(FM_L5L6_L1_FromMinus_FT_L5L6_read_en),
.fullmatch1in4(FM_L5L6_L1_FromMinus_FT_L5L6),
.number2in4(FM_L5L6_L2_FromMinus_FT_L5L6_number),
.read_add2in4(FM_L5L6_L2_FromMinus_FT_L5L6_read_add),
.read_en2in4(FM_L5L6_L2_FromMinus_FT_L5L6_read_en),
.fullmatch2in4(FM_L5L6_L2_FromMinus_FT_L5L6),
.number3in4(FM_L5L6_L3_FromMinus_FT_L5L6_number),
.read_add3in4(FM_L5L6_L3_FromMinus_FT_L5L6_read_add),
.read_en3in4(FM_L5L6_L3_FromMinus_FT_L5L6_read_en),
.fullmatch3in4(FM_L5L6_L3_FromMinus_FT_L5L6),
.number4in4(FM_L5L6_L4_FromMinus_FT_L5L6_number),
.read_add4in4(FM_L5L6_L4_FromMinus_FT_L5L6_read_add),
.read_en4in4(FM_L5L6_L4_FromMinus_FT_L5L6_read_en),
.fullmatch4in4(FM_L5L6_L4_FromMinus_FT_L5L6),
.trackout(FT_L5L6_TF_L5L6),
.valid_fit(FT_L5L6_TF_L5L6_wr_en),
.start(FM_L5L6_L4_FromMinus_start),
.done(FT_L5L6_start),
.clk(clk),
.clk_new(clk_new),		  //MT			   
.reset(reset),
.en_proc(en_proc)
);

PurgeDuplicate #(.SCOPE("D3D4")) PD(
.numberin1(TF_L1L2_PD_number),
.read_add_trackin1(TF_L1L2_PD_read_add),
.index_in1(TF_L1L2_PD_index),
.trackin1(TF_L1L2_PD),
.numberin2(TF_L3L4_PD_number),
.read_add_trackin2(TF_L3L4_PD_read_add),
.index_in2(TF_L3L4_PD_index),
.trackin2(TF_L3L4_PD),
.numberin3(TF_L5L6_PD_number),
.read_add_trackin3(TF_L5L6_PD_read_add),
.index_in3(TF_L5L6_PD_index),
.trackin3(TF_L5L6_PD),
.trackout1(PD_CT_L1L2),
.trackout2(PD_CT_L3L4),
.trackout3(PD_CT_L5L6),
.valid_out_1(PD_CT_L1L2_wr_en),
.valid_out_2(PD_CT_L3L4_wr_en),
.valid_out_3(PD_CT_L5L6_wr_en),
.start(TF_L1L2_start),
.done(PD_start),
.clk(clk),
.reset(reset),
.en_proc(en_proc)
);

wire [31:0] reader_out;

wire InputLink_R1Link1_io_rd_ack , InputLink_R1Link2_io_rd_ack , InputLink_R1Link3_io_rd_ack;
wire TPars_L1L2_io_rd_ack , TPars_L3L4_io_rd_ack , TPars_L5L6_io_rd_ack;
// readback mux
// If a particular block is addressed, connect that block's signals
// to the 'rdbk' output. At the same time, assert 'rdbk_sel' to tell downstream muxes to
// use the 'rdbk' from this module as their source of data.
reg [31:0] io_rd_data_reg;
assign io_rd_data = io_rd_data_reg;
// Assert 'io_rd_ack' if any module is asserting its 'rd_ack'.
reg io_rd_ack_reg;
assign io_rd_ack = io_rd_ack_reg;
always @ (posedge io_clk) begin
io_rd_ack_reg <= InputLink_R1Link1_io_rd_ack | InputLink_R1Link2_io_rd_ack | InputLink_R1Link3_io_rd_ack |
TPars_L1L2_io_rd_ack | TPars_L3L4_io_rd_ack | TPars_L5L6_io_rd_ack;
end
// Route the selected register to the 'rdbk' output.
always @(posedge io_clk) begin
if (InputLink_R1Link1_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link1_io_rd_data[31:0];
if (InputLink_R1Link2_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link2_io_rd_data[31:0];
if (InputLink_R1Link3_io_sel) io_rd_data_reg[31:0] <= InputLink_R1Link3_io_rd_data[31:0];
if (TPars_L1L2_io_sel) io_rd_data_reg[31:0] <= TPars_L1L2_io_rd_data[31:0];
if (TPars_L3L4_io_sel) io_rd_data_reg[31:0] <= TPars_L3L4_io_rd_data[31:0];
if (TPars_L5L6_io_sel) io_rd_data_reg[31:0] <= TPars_L5L6_io_rd_data[31:0];
//if (reader_ack)    io_rd_data_reg <= reader_out;
end

endmodule
